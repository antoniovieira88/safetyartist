library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 0, 2, 1, 0, 1, 0, -2, -2, -2, 1, -2, 1, -2, 1, -2, -2, 1, 0, -2, 0, 1, -2, -2, 0, -2, -2, 1, 0, -2, -2, -2, 2, 0, 0, 0, -2, 1, -2, -2, 1, 1, -2, -2, 1, -2, -2, 0, 1, 0, -2, -2, 1, -2, -2, -2, 0, 0, 0, 0, -2, -2, 0, -2, -2, 1, -2, 1, -2, -2, 0, 0, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, 1, -2, -2, 2, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, 1, -2, 0, 1, -2, 1, -2, -2, -2, 2, 1, 1, -2, 0, -2, -2, 0, 1, 1, -2, -2, -2, 0, 1, -2, -2, -2, 1, 0, 1, -2, -2, -2, 0, 1, 1, -2, -2, -2, -2, 0, 2, 1, 0, 0, -2, 0, -2, 1, -2, -2, 1, 1, -2, 1, -2, -2, 0, -2, 1, -2, -2, 1, 0, -2, -2, -2, 0, 1, 0, 1, 0, -2, -2, 1, -2, -2, -2, -2, 0, 1, 0, 1, -2, -2, 0, -2, -2, -2, 1, -2, -2, 2, 1, 0, 1, -2, 0, -2, 1, -2, -2, -2, 1, -2, 1, 0, -2, -2, 1, -2, 0, -2, -2, 1, 0, 0, -2, -2, -2, 0, 0, -2, 1, -2, -2, 1, -2, 1, 0, -2, -2, -2, 2, 0, 2, 0, 0, 0, -2, 1, -2, -2, 0, -2, 0, -2, 1, -2, -2, 1, 1, -2, 1, -2, 0, -2, -2, 0, 0, -2, 0, -2, -2, 1, 0, -2, -2, -2, 2, 1, 0, 1, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, -2, 1, 1, 0, -2, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 1, 0, -2, 0, -2, -2, -2, 1, 1, -2, 1, -2, -2, 1, 1, -2, -2, 1, -2, -2, 0, 1, 2, 0, 1, -2, 0, -2, -2, 1, -2, 0, -2, -2, -2, 0, 1, 0, 0, -2, -2, -2, 0, 0, -2, -2, 2, -2, -2, 1, 1, 2, -2, -2, 1, -2, -2, 1, 1, -2, -2, -2, 1, 1, -2, 0, 2, 1, -2, -2, 0, -2, -2, 1, -2, 2, -2, -2, 2, 1, 1, -2, 0, -2, -2, 1, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, -2, 1, 0, 2, 1, 1, 0, -2, -2, -2, 1, 0, -2, -2, 1, 0, -2, -2, -2, 0, 1, 0, -2, -2, 1, 0, -2, -2, -2, 0, 0, 1, -2, -2, -2, 0, -2, 0, -2, -2, 1, 2, 0, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, 1, 1, -2, 1, -2, -2, 1, -2, -2, 2, 0, -2, -2, 0, -2, 1, -2, 0, -2, -2, 2, 1, 0, -2, -2, 1, 1, 0, 0, -2, -2, 1, -2, -2, 0, -2, -2, 1, -2, 0, -2, -2, 0, 0, -2, 1, 1, 1, -2, -2, -2, -2, 1, -2, 1, -2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 0, 1, 1, 0, 1, 2, 1, 0, -2, -2, -2, 0, -2, -2, 2, 1, 1, -2, -2, -2, 0, -2, 1, -2, -2, 2, 1, 1, -2, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, -2, 0, 2, 1, 1, 1, -2, -2, -2, -2, 0, -2, 1, 0, -2, -2, -2, 0, 1, 2, 0, -2, -2, -2, 1, 1, -2, -2, -2, 2, 0, 0, -2, -2, -2, -2, 2, 0, 0, -2, 0, -2, 0, 1, -2, -2, 0, -2, -2, 0, 0, 1, 0, -2, -2, -2, -2, 0, -2, 1, -2, -2, 1, 0, 1, 1, -2, -2, -2, 1, 0, 0, -2, -2, -2, 1, 0, -2, -2, 1, -2, -2, 0, -2, 0, -2, 1, -2, 1, -2, -2, 0, 1, 2, 1, 1, 1, -2, 1, -2, -2, 1, -2, 1, -2, -2, 1, 0, 1, -2, -2, 0, -2, -2, 0, -2, -2, 1, 1, -2, 0, -2, -2, 1, 0, 1, -2, -2, 1, -2, -2, 1, -2, 1, -2, -2, 1, 0, -2, 0, -2, 0, 1, -2, -2, -2, 2, -2, 1, 1, -2, 1, -2, -2, 1, 1, -2, -2, -2, 1, 2, 1, 0, 0, -2, -2, -2, 1, -2, 1, 0, -2, -2, 1, -2, -2, -2, 1, -2, 0, 2, 1, 1, -2, -2, 0, -2, -2, 0, 0, -2, -2, -2, -2, 1, 1, 1, 1, 0, 2, 0, -2, 0, -2, -2, 0, -2, 0, -2, -2, 1, -2, 1, -2, 1, -2, -2, 2, 1, 1, 0, -2, -2, -2, 1, -2, 1, -2, -2, 2, 0, -2, -2, 1, -2, 1, -2, -2, 0, 2, 0, -2, 1, -2, -2, 2, 1, 0, -2, -2, -2, 0, -2, 0, -2, -2, 1, 0, 1, -2, 1, -2, -2, -2, 2, 1, -2, 0, -2, -2, 0, -2, 1, -2, -2, 1, -2, 0, 2, 1, 1, -2, 0, -2, -2, -2, 1, 1, 2, -2, -2, 2, -2, -2, 2, -2, 0, -2, -2, 0, 0, 2, 0, -2, -2, 1, -2, -2, 0, 0, -2, -2, -2, 1, 1, -2, 1, -2, -2, 1, 0, -2, -2, 0, -2, -2, 1, 0, 2, -2, 1, 0, 2, -2, 1, -2, -2, 1, 1, -2, -2, -2, 1, 1, 2, -2, -2, -2, 0, 0, -2, -2, 2, -2, -2, 2, 1, 0, 1, 0, -2, -2, -2, 1, 1, -2, -2, -2, 1, -2, 1, 0, -2, -2, 1, -2, -2, 2, 0, 1, -2, 1, -2, -2, -2, -2, 1, 1, 2, 2, 0, -2, -2, 1, -2, -2, 1, -2, -2, 2, 2, 0, 1, -2, -2, 1, -2, -2, 1, 0, -2, -2, 0, -2, -2, 0, 0, -2, 0, -2, -2, 1, 0, -2, -2, 0, -2, -2, 2, 0, 1, 1, 1, -2, -2, -2, 0, -2, -2, -2, 0, 0, 0, -2, 2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 1, 2, 0, 0, 0, -2, 0, 0, -2, -2, 1, -2, -2, 1, -2, -2, 0, 1, 1, -2, 1, -2, -2, 0, -2, 1, -2, -2, 1, -2, 0, -2, -2, 2, 1, 0, 1, 0, -2, -2, 0, -2, -2, -2, 0, 0, -2, 1, -2, -2, 1, -2, 1, -2, -2, 0, 1, 1, 0, -2, -2, -2, 1, 1, -2, -2, -2, 0, 1, 0, -2, -2, 0, -2, -2, -2, 1, 1, 0, -2, -2, 2, 1, 1, 1, -2, -2, -2, 1, 0, -2, -2, 0, -2, -2, 2, 1, 0, -2, -2, -2, 0, 0, -2, -2, 1, -2, -2, 1, -2, 2, 0, 0, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, 0, -2, -2, 2, 1, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 0, 2, 0, -2, 0, -2, 1, -2, 0, -2, -2, 1, 1, 1, 0, -2, -2, -2, 0, -2, -2, -2, 1, 1, 0, 2, 1, -2, -2, -2, -2, 1, -2, 0, -2, 0, -2, -2, 1, 0, 0, -2, 2, -2, -2, -2, -2, 2, 1, 1, -2, 1, -2, 1, 1, -2, -2, 0, -2, -2, 1, -2, 1, 1, 1, -2, -2, 0, -2, -2, 1, -2, 1, -2, -2, 1, 1, 1, -2, 1, -2, -2, 0, 1, 1, -2, -2, -2, -2, 1, -2, 1, 0, -2, -2, -2, 2, 1, 0, 0, 1, 1, 1, 2, -2, -2, 1, -2, -2, -2, 1, 0, -2, 0, -2, -2, -2, 1, 2, 1, -2, 1, -2, -2, -2, 0, 2, -2, 1, -2, -2, 2, -2, 0, -2, -2, 1, -2, 1, 0, -2, -2, 1, 0, 2, -2, -2, -2, 2, 1, -2, -2, -2, 2, 1, 1, 1, 0, 1, -2, -2, -2, -2, 1, 0, -2, -2, 0, 0, -2, -2, 0, -2, -2, 1, 1, -2, 0, -2, -2, 1, -2, 1, 1, -2, -2, 1, -2, -2, 1, 1, 1, 0, 1, -2, -2, 0, -2, -2, 1, -2, 0, -2, -2, 1, 1, 0, -2, -2, -2, 0, -2, -2, 1, 0, -2, -2, -2, 2, 1, 0, -2, 1, 0, 0, -2, 0, -2, -2, -2, 1, -2, 0, -2, -2, 1, 1, 1, 0, -2, -2, 1, 0, -2, -2, 1, -2, -2, 0, 0, 0, -2, -2, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, 1, -2, 1, 1, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 2, 1, -2, 0, 1, 0, 0, -2, -2, 0, -2, -2, 1, 1, -2, -2, 0, -2, -2, 1, -2, 1, -2, 1, -2, -2, 1, 0, 1, 1, -2, -2, -2, -2, 0, 1, 0, 0, -2, -2, 1, -2, -2, -2, 1, 0, 0, -2, -2, -2, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((2202, 134, 19321, 92, 1021, 3973, 449, 1247, -256, -256, -256, 644, -256, 665, -256, 918, -256, -256, 1372, 11695, -256, 13014, 1144, -256, -256, 15847, -256, -256, 1439, 15958, -256, -256, -256, 109, 8073, 2377, 1118, -256, 337, -256, -256, 734, 506, -256, -256, 930, -256, -256, 19255, 1396, 13437, -256, -256, 1607, -256, -256, -256, 7553, 3701, 2427, 1179, -256, -256, 2433, -256, -256, 708, -256, 886, -256, -256, 12829, 7808, 993, -256, -256, 1086, -256, -256, 14184, 13769, -256, -256, 1582, -256, -256, 92, 29241, 29143, 28076, 27884, 26723, -256, -256, -256, -256, -256, 2045, -256, 34655, 2048, -256, 2078, -256, -256, -256, 109, 1890, 1740, -256, 22444, -256, -256, 27433, 1934, 1901, -256, -256, -256, 30086, 2031, -256, -256, -256, 1880, 20294, 1754, -256, -256, -256, 26887, 2084, 2068, -256, -256, -256, -256, 12732, 164, 1132, 3726, 1348, -256, 1359, -256, 361, -256, -256, 810, 608, -256, 618, -256, -256, 6435, -256, 1025, -256, -256, 1333, 10891, -256, -256, -256, 4968, 687, 2501, 33, 626, -256, -256, 329, -256, -256, -256, -256, 11424, 1208, 6158, 864, -256, -256, 7701, -256, -256, -256, 1555, -256, -256, 164, 1937, 18098, 1628, -256, 16049, -256, 1793, -256, -256, -256, 1937, -256, 2004, 21208, -256, -256, 2005, -256, 23085, -256, -256, 1771, 13522, 13163, -256, -256, -256, 19162, 15968, -256, 1942, -256, -256, 2045, -256, 2046, 136555, -256, -256, -256, 134, 57867, 92, 42531, 39695, 37207, -256, 2221, -256, -256, 39730, -256, 42284, -256, 2548, -256, -256, 2748, 2498, -256, 2514, -256, 52390, -256, -256, 57440, 55098, -256, 55167, -256, -256, 2964, 57646, -256, -256, -256, 109, 2641, 40059, 2228, 2227, -256, -256, 37775, -256, -256, 42127, 2489, -256, -256, -256, 2835, 2835, 47368, -256, -256, -256, 54836, 2874, -256, -256, 3059, -256, -256, 35932, 2402, 29842, -256, 32751, -256, -256, -256, 2787, 2593, -256, 2615, -256, -256, 3002, 2964, -256, -256, 3314, -256, -256, 73034, 3068, 92, 62717, 2798, -256, 59422, -256, -256, 3047, -256, 70409, -256, -256, -256, 64473, 3141, 59718, 58389, -256, -256, -256, 63885, 62540, -256, -256, 109, -256, -256, 3529, 3164, 92, -256, -256, 3287, -256, -256, 3713, 3562, -256, -256, -256, 3411, 3247, -256, 78000, 92, 3319, -256, -256, 75662, -256, -256, 3248, -256, 92, -256, -256, 92, 3413, 3412, -256, 119687, -256, -256, 3789, 86465, -256, -256, 116240, -256, -256, 74093, 3466, -256, -256, -256, 3085, 31814, 164, 2314, 2311, 26368, -256, -256, -256, 2442, 28216, -256, -256, 2576, 29493, -256, -256, -256, 26660, 2230, 22490, -256, -256, 2495, 24009, -256, -256, -256, 30750, 30614, 2664, -256, -256, -256, 31297, -256, 31762, -256, -256, 2884, 164, 33391, 2566, -256, -256, 2791, 34743, -256, -256, 2792, -256, -256, 2871, 2744, -256, 2745, -256, -256, 2871, -256, -256, 164, 41057, -256, -256, 35977, -256, 3040, -256, 41619, -256, -256, 164, 3125, 43933, -256, -256, 3680, 3668, 52715, 50994, -256, -256, 3461, -256, -256, 69086, -256, -256, 3729, -256, 57374, -256, -256, 44762, 40818, -256, 3339, 3250, 3167, -256, -256, -256, -256, 3455, -256, 3456, -256, 48162, 3497, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256),
                (109, 42413, 1693, 928, 3869, 270, 92, 264, 1247, -256, -256, -256, 1159, -256, -256, 92, 541, 506, -256, -256, -256, 1937, -256, 489, -256, -256, 92, 918, 646, -256, 5789, -256, -256, 20432, -256, -256, 4881, 668, -256, -256, -256, 15438, 92, 1264, 1257, 1065, -256, -256, -256, -256, 9881, -256, 1287, 12271, -256, -256, -256, 19308, 1443, 92, 16714, -256, -256, -256, 1538, 1526, -256, -256, -256, 92, 24250, 24108, -256, -256, -256, -256, 92, 31972, 26752, -256, 26774, -256, 30441, 1919, -256, -256, 31852, -256, -256, 42309, 42135, 2222, 35249, -256, -256, -256, -256, 42360, -256, 2290, -256, -256, 2215, 25078, 1733, 1729, -256, -256, -256, 2026, 26772, 26712, -256, -256, -256, 2065, 33308, -256, -256, 2110, -256, -256, 37250, -256, 37319, -256, 2412, -256, 2588, -256, -256, 71826, 3006, 92, 2724, 2465, 2371, -256, 2383, -256, -256, 2471, -256, 2676, -256, -256, 2956, 60676, 2873, -256, -256, 62166, -256, -256, 61451, -256, -256, 2808, 2730, -256, 46635, -256, -256, 2870, 53696, 2834, -256, -256, 2831, -256, -256, 2891, -256, 2897, -256, -256, 3066, 63263, -256, 66580, -256, 69250, 3024, -256, -256, -256, 92, -256, 3417, 3084, -256, 3331, -256, -256, 3491, 3479, -256, -256, -256, 3404, 92, 3280, 75496, 75491, -256, -256, -256, 3281, -256, 3307, 80659, -256, -256, 3361, -256, -256, -256, 3404, -256, 89603, 92, 3438, 3424, -256, -256, 87034, -256, -256, 72928, 72733, -256, -256, -256, -256, 2402, 1643, 906, 516, 2455, 134, 1297, -256, 1362, -256, -256, 1142, -256, 1263, -256, -256, 441, -256, 441, -256, 451, -256, -256, 134, 842, 842, 5200, -256, -256, -256, 890, -256, 890, -256, -256, 164, 3903, -256, -256, 516, -256, 570, -256, -256, 9519, 134, 8906, -256, 1229, -256, -256, 164, 1093, 6901, -256, -256, -256, 6507, -256, 7471, -256, -256, 1343, 11453, 1229, -256, 1303, -256, -256, -256, 164, 1343, -256, 13294, -256, -256, 10930, -256, 1457, -256, -256, 1643, -256, 21001, 134, 1664, 1652, -256, 14600, -256, -256, -256, 1982, 1973, 164, -256, -256, 164, -256, -256, 164, -256, 17202, -256, -256, 24550, 21782, 134, 21725, -256, -256, 2146, -256, -256, 24399, 23126, -256, -256, -256, 2166, 2056, -256, 2056, -256, -256, 2172, 27460, -256, -256, 29449, -256, -256, 2884, 34494, 134, -256, 2595, 28721, 164, -256, 2595, -256, -256, 2539, 2493, -256, -256, -256, 2676, 2673, 164, -256, -256, -256, 34304, 32014, -256, -256, 164, -256, -256, 134, 2798, 37616, 2603, 36003, -256, -256, -256, 2593, 2592, -256, -256, -256, 2798, -256, 2799, 42104, -256, -256, 2873, -256, -256, 164, 38090, 2667, -256, 2864, -256, -256, -256, -256, 3474, 2887, 164, 134, 60789, -256, -256, 2886, -256, -256, 2886, -256, -256, 164, 134, 55642, 2894, -256, -256, 3462, -256, -256, 2901, 44890, -256, -256, 48339, -256, -256, 40855, 35943, -256, 36126, -256, -256, 3430, 42312, -256, -256, 46871, -256, -256, 134, 66423, 3648, 3502, 3499, -256, -256, -256, 61338, -256, -256, -256, 54447, 48741, 46034, -256, 164, -256, -256, 164, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256),
                (2362, 134, 1357, 92, 5255, 3635, 1269, -256, 1321, 1310, -256, -256, 339, -256, -256, 569, -256, -256, 11695, 920, 744, -256, 807, -256, -256, 10227, -256, 1023, -256, -256, 1228, -256, 14501, -256, -256, 109, 926, 4881, 538, 1116, -256, -256, 4723, -256, -256, -256, 9612, 8330, -256, 1013, -256, -256, 1224, -256, 1226, -256, -256, 5314, 434, 383, 693, -256, -256, -256, 686, 671, -256, -256, -256, 11419, 1001, 7833, -256, -256, 10130, -256, -256, -256, 1916, 1358, 81991, -256, -256, 92, 1880, 1879, 1544, -256, -256, -256, 1914, 20726, -256, -256, 28479, -256, -256, 109, 1893, 18990, -256, -256, -256, 15972, 14165, -256, -256, 1744, -256, -256, 1916, -256, 92, 35806, 33120, 1952, -256, -256, 2113, -256, -256, 38932, 38303, -256, -256, 44761, -256, -256, 109, 2079, 1949, -256, -256, 30966, -256, -256, 26872, 2080, -256, -256, 2319, -256, -256, 12899, 3691, 164, 1243, -256, 1248, -256, 226, -256, 2640, -256, -256, 255, 67, 64, 1255, -256, -256, -256, 612, -256, -256, -256, 1225, 843, 4930, 164, 608, -256, -256, -256, -256, 844, -256, 6322, -256, 8263, -256, -256, 1383, 11279, 9557, -256, 164, -256, -256, -256, -256, 164, 1915, 1638, -256, 1639, -256, 1724, 1724, -256, -256, 17222, -256, -256, 1915, -256, 2248, 1923, 1922, -256, -256, 21872, -256, -256, 2249, -256, 2250, -256, -256, 2203, 1807, 1567, -256, 1568, -256, -256, 19075, 1882, 1855, -256, -256, -256, -256, 2205, -256, 2336, 23122, -256, -256, -256, 109, 3028, 52307, 45839, 2468, 2467, 2391, 92, -256, -256, 2392, -256, -256, -256, 2625, 42642, -256, 43371, -256, -256, -256, 2610, 92, 2440, -256, 2559, -256, -256, -256, 48791, 92, -256, 2818, -256, -256, 92, -256, 49472, -256, -256, 2767, -256, 2768, 97902, -256, -256, 2906, 62717, 92, -256, -256, -256, 92, 2961, -256, -256, -256, 92, 3556, 3052, 3052, 69099, 3042, -256, -256, -256, -256, 3128, 71567, -256, -256, 75724, 74128, -256, -256, 81958, -256, -256, 3577, 3561, -256, 85867, -256, -256, 3584, -256, 3685, 3677, -256, -256, 3698, -256, -256, 3657, 3582, 3578, 67955, 3091, -256, -256, 73025, -256, -256, 3579, -256, 84053, -256, -256, 3618, 3601, 69362, -256, -256, -256, 67314, -256, -256, 3734, 75593, -256, -256, -256, 134, 2665, 33403, -256, 2437, 36658, 33925, -256, 36006, -256, -256, -256, 2593, -256, 39895, -256, -256, 3250, 2694, 2689, 39078, -256, -256, 2692, 91368, -256, -256, 2693, -256, -256, 47238, 44067, 43445, -256, -256, 2817, -256, -256, 3039, 51306, -256, -256, 3040, -256, -256, 3250, -256, 3281, 3260, 57582, -256, -256, 59525, -256, -256, 63956, 3284, -256, -256, 65327, -256, -256, 164, 2363, -256, 43495, 2663, 30177, 28943, -256, -256, 30644, -256, -256, 2805, 2792, -256, -256, 41048, -256, -256, 3185, -256, 3186, -256, 3187, -256, -256, 2616, 27370, 2377, 2375, -256, -256, -256, -256, 40855, 3076, 33107, 30633, -256, -256, 2882, -256, -256, -256, 3429, 42371, 42262, -256, -256, -256, 3429, -256, 3439, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((38, 41, 41, 19, 18, 34, 9, 22, 0, 43, 0, 40, 43, 34, 0, 35, 37, 30, 4, 13, 0, 37, 21, 43, 0, 40, 35, 43, 0, 4, 0, 43, 0, 19, 19, 11, 2, 0, 4, 43, 0, 14, 38, 43, 24, 2, 14, 0, 26, 26, 39, 35, 42, 2, 6, 0, 0, 18, 9, 3, 1, 0, 3, 7, 43, 5, 15, 43, 2, 13, 0, 25, 21, 32, 43, 0, 19, 41, 1, 28, 36, 29, 41, 26, 42, 1, 42, 42, 32, 33, 32, 32, 32, 38, 0, 43, 0, 43, 43, 42, 6, 0, 11, 43, 0, 43, 42, 42, 43, 43, 42, 0, 43, 41, 5, 21, 0, 43, 0, 43, 30, 43, 0, 43, 43, 43, 41, 43, 0, 43, 42, 5, 9, 4, 43, 0, 43, 41, 17, 17, 29, 6, 0, 13, 43, 11, 43, 0, 37, 41, 43, 38, 0, 41, 27, 0, 41, 43, 39, 1, 7, 0, 43, 0, 17, 6, 19, 6, 28, 0, 43, 3, 9, 0, 43, 0, 24, 22, 40, 34, 43, 0, 42, 41, 43, 0, 31, 43, 0, 42, 42, 43, 40, 43, 12, 0, 26, 43, 0, 43, 41, 0, 41, 42, 0, 43, 40, 0, 41, 0, 43, 42, 43, 41, 43, 0, 43, 42, 5, 0, 14, 43, 0, 43, 43, 43, 32, 0, 43, 43, 34, 33, 6, 4, 0, 0, 0, 1, 43, 0, 3, 43, 1, 0, 6, 43, 0, 15, 37, 43, 28, 0, 31, 13, 43, 1, 0, 0, 2, 43, 0, 9, 16, 43, 0, 0, 7, 6, 16, 2, 20, 16, 43, 1, 0, 9, 40, 27, 43, 0, 43, 2, 6, 6, 0, 39, 43, 1, 0, 1, 0, 7, 38, 0, 7, 0, 3, 0, 32, 21, 43, 0, 20, 40, 43, 36, 14, 37, 7, 18, 15, 43, 4, 6, 0, 42, 31, 41, 39, 28, 43, 3, 21, 0, 42, 43, 32, 0, 43, 43, 14, 7, 35, 28, 43, 0, 43, 4, 3, 5, 0, 11, 0, 32, 21, 24, 13, 3, 43, 27, 39, 21, 8, 7, 0, 9, 43, 42, 43, 43, 42, 29, 6, 0, 14, 40, 43, 32, 43, 0, 43, 43, 43, 42, 39, 14, 0, 21, 0, 43, 40, 40, 2, 43, 27, 0, 43, 43, 28, 0, 43, 43, 36, 37, 3, 1, 7, 6, 0, 43, 43, 0, 2, 0, 43, 0, 1, 0, 9, 0, 4, 1, 6, 0, 43, 0, 2, 0, 26, 0, 22, 27, 25, 41, 0, 43, 4, 0, 14, 43, 0, 42, 43, 42, 21, 43, 0, 43, 43, 37, 43, 42, 0, 42, 43, 43, 43, 42, 0, 43, 42, 0, 43, 42, 41, 0, 43, 42, 0, 43, 43, 42, 21, 43, 34, 34, 28, 0, 43, 34, 34, 34, 1, 0, 20, 43, 43, 42, 16, 0, 43, 42, 43, 39, 0, 43, 35, 1, 0, 15, 38, 34, 43, 0, 43, 0, 43, 43, 42, 0, 42, 21, 43, 14, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43),
                (38, 38, 18, 34, 39, 12, 29, 32, 30, 0, 43, 43, 25, 0, 43, 4, 4, 9, 4, 43, 0, 4, 0, 11, 43, 0, 42, 42, 42, 43, 41, 0, 42, 21, 0, 43, 42, 28, 43, 0, 43, 28, 6, 5, 10, 9, 5, 12, 43, 0, 7, 0, 18, 38, 30, 43, 0, 41, 32, 41, 39, 26, 43, 43, 3, 11, 0, 43, 0, 42, 42, 39, 40, 0, 43, 43, 4, 3, 1, 0, 4, 43, 4, 5, 43, 0, 1, 0, 4, 11, 10, 11, 36, 24, 43, 0, 0, 21, 43, 16, 43, 0, 4, 14, 0, 7, 0, 43, 0, 38, 41, 32, 37, 0, 43, 30, 14, 0, 43, 37, 43, 34, 1, 0, 6, 43, 5, 43, 1, 7, 0, 41, 34, 41, 40, 42, 43, 43, 41, 0, 43, 33, 0, 34, 32, 43, 18, 16, 3, 4, 0, 39, 26, 43, 31, 0, 43, 41, 43, 43, 36, 0, 43, 28, 19, 3, 21, 0, 39, 32, 43, 31, 43, 29, 0, 32, 4, 19, 0, 35, 43, 24, 11, 43, 0, 43, 2, 0, 5, 9, 43, 8, 6, 16, 1, 1, 0, 43, 0, 43, 43, 43, 43, 42, 43, 0, 43, 41, 0, 41, 40, 0, 43, 42, 42, 43, 43, 41, 0, 41, 24, 2, 14, 0, 43, 1, 0, 9, 40, 24, 43, 0, 43, 43, 39, 41, 42, 42, 42, 7, 6, 0, 21, 43, 14, 8, 0, 24, 43, 0, 43, 43, 43, 0, 43, 42, 43, 42, 42, 42, 42, 2, 43, 0, 42, 43, 42, 0, 43, 42, 42, 0, 43, 42, 0, 42, 40, 42, 41, 3, 0, 0, 11, 43, 0, 4, 5, 16, 0, 43, 0, 3, 0, 20, 43, 12, 42, 43, 37, 43, 9, 0, 43, 43, 42, 42, 0, 42, 0, 43, 42, 0, 43, 43, 43, 39, 0, 39, 3, 0, 11, 0, 28, 0, 43, 0, 4, 8, 7, 7, 8, 32, 0, 43, 0, 0, 1, 0, 3, 42, 25, 36, 38, 43, 0, 34, 43, 0, 22, 23, 17, 28, 0, 43, 43, 43, 43, 0, 43, 42, 41, 17, 43, 42, 30, 43, 35, 37, 4, 0, 5, 10, 2, 0, 5, 3, 43, 39, 37, 43, 21, 43, 2, 4, 1, 0, 1, 43, 1, 0, 0, 5, 21, 0, 43, 42, 42, 42, 15, 27, 43, 17, 0, 43, 42, 43, 0, 43, 40, 0, 41, 32, 0, 43, 41, 40, 43, 43, 42, 33, 43, 19, 14, 43, 43, 43, 34, 35, 19, 17, 17, 0, 43, 17, 0, 43, 21, 43, 0, 35, 34, 34, 2, 21, 2, 42, 42, 37, 35, 39, 0, 43, 34, 2, 43, 36, 2, 0, 17, 43, 14, 42, 43, 30, 43, 40, 14, 43, 32, 31, 1, 0, 2, 0, 43, 0, 5, 0, 43, 43, 33, 2, 0, 0, 7, 0, 21, 16, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
                (39, 41, 40, 42, 42, 10, 4, 0, 8, 28, 43, 21, 5, 43, 0, 19, 43, 0, 42, 30, 42, 43, 35, 14, 43, 1, 0, 6, 43, 0, 43, 43, 42, 0, 43, 42, 42, 42, 17, 28, 0, 40, 2, 0, 14, 43, 41, 1, 0, 14, 43, 0, 42, 43, 42, 0, 42, 42, 11, 28, 25, 0, 41, 43, 2, 8, 6, 43, 0, 42, 31, 41, 40, 43, 4, 0, 21, 43, 39, 39, 9, 0, 43, 39, 39, 39, 39, 40, 38, 0, 42, 42, 0, 43, 38, 0, 43, 40, 40, 39, 1, 42, 43, 40, 2, 0, 12, 42, 43, 42, 38, 0, 38, 37, 2, 0, 2, 0, 18, 43, 0, 42, 30, 36, 18, 43, 41, 43, 38, 38, 39, 37, 40, 37, 0, 42, 38, 0, 1, 0, 42, 43, 41, 41, 15, 3, 3, 0, 5, 43, 5, 43, 1, 0, 3, 3, 26, 14, 28, 0, 43, 0, 33, 0, 43, 0, 20, 37, 42, 37, 33, 43, 0, 43, 43, 28, 0, 29, 0, 38, 28, 43, 2, 16, 2, 0, 11, 0, 43, 43, 0, 42, 42, 43, 43, 42, 0, 42, 42, 42, 0, 42, 0, 43, 41, 0, 41, 41, 37, 43, 0, 42, 0, 43, 40, 0, 40, 36, 40, 42, 43, 43, 43, 43, 0, 43, 42, 6, 16, 7, 43, 0, 43, 41, 0, 41, 40, 0, 43, 43, 34, 33, 34, 3, 1, 3, 2, 1, 0, 3, 3, 43, 2, 43, 0, 0, 0, 12, 43, 7, 0, 19, 35, 28, 43, 18, 0, 43, 43, 8, 14, 0, 30, 36, 0, 3, 0, 14, 0, 17, 42, 43, 42, 28, 0, 43, 42, 41, 23, 15, 36, 43, 42, 42, 42, 42, 43, 31, 30, 31, 25, 26, 1, 3, 0, 43, 0, 31, 33, 0, 43, 30, 0, 0, 7, 42, 29, 42, 24, 8, 0, 12, 0, 43, 26, 43, 25, 23, 24, 0, 31, 43, 26, 32, 33, 32, 33, 3, 11, 1, 42, 30, 43, 16, 0, 21, 0, 43, 37, 41, 40, 0, 43, 43, 32, 0, 43, 25, 22, 0, 43, 43, 36, 35, 37, 0, 42, 42, 21, 43, 11, 21, 0, 43, 42, 43, 42, 0, 43, 34, 34, 30, 33, 0, 43, 15, 7, 0, 43, 21, 43, 14, 35, 1, 0, 0, 5, 17, 43, 7, 42, 43, 39, 43, 42, 0, 42, 32, 0, 33, 28, 37, 0, 43, 21, 0, 43, 33, 2, 43, 2, 43, 24, 43, 36, 36, 0, 36, 5, 13, 0, 0, 11, 41, 21, 42, 1, 6, 4, 17, 1, 0, 9, 42, 43, 41, 0, 42, 32, 42, 37, 39, 1, 9, 0, 43, 0, 43, 36, 3, 7, 1, 0, 11, 35, 43, 26, 0, 42, 43, 33, 38, 0, 43, 42, 0, 42, 39, 42, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 3, 4, 5, 6, 7, 8, 505, 507, 509, 12, 511, 14, 513, 16, -1, -1, 19, 20, 515, 22, 23, -1, -1, 26, -1, -1, 29, 30, 517, 519, 521, 34, 35, 36, 37, 523, 39, -1, -1, 42, 43, -1, -1, 46, -1, -1, 49, 50, 51, -1, -1, 54, -1, -1, 525, 58, 59, 60, 61, -1, -1, 64, -1, -1, 67, 527, 69, -1, -1, 72, 73, 74, -1, -1, 77, -1, -1, 80, 81, -1, -1, 84, -1, -1, 87, 88, 89, 90, 91, 92, -1, -1, 529, 531, 533, 98, 535, 100, 101, 537, 103, -1, -1, 539, 107, 108, 109, 541, 111, 543, 545, 114, 115, 116, -1, -1, 547, 120, 121, -1, -1, 549, 125, 126, 127, 551, 553, 555, 131, 132, 133, -1, -1, 557, 559, 138, 139, 140, 141, 142, 561, 144, 563, 146, -1, -1, 149, 150, 565, 152, -1, -1, 155, 567, 157, -1, -1, 160, 161, 569, 571, 573, 165, 166, 167, 168, 169, -1, -1, 172, -1, -1, 575, 577, 177, 178, 179, 180, -1, -1, 183, -1, -1, 579, 187, 581, 583, 190, 191, 192, 193, 585, 195, 587, 197, -1, -1, 589, 201, 591, 203, 204, 593, 595, 207, 597, 209, -1, -1, 212, 213, 214, 599, 601, 603, 218, 219, 605, 221, 607, 609, 224, 611, 226, 227, -1, -1, 613, 231, 232, 233, 234, 235, 236, 615, 238, 617, 619, 241, 621, 243, 623, 245, -1, -1, 248, 249, 625, 251, 627, 253, -1, -1, 256, 257, 629, 259, -1, -1, 262, 263, -1, -1, 631, 267, 268, 269, 270, 271, -1, -1, 274, -1, -1, 277, 278, -1, -1, 633, 282, 283, 284, -1, -1, 635, 288, 289, -1, -1, 292, -1, -1, 295, 296, 297, 637, 299, -1, -1, 639, 303, 304, 641, 306, -1, -1, 309, 310, -1, -1, 313, -1, -1, 316, 317, 318, 319, 320, 643, 322, -1, -1, 325, 645, 327, -1, -1, 647, 331, 332, 333, 334, -1, -1, 649, 338, 339, -1, -1, 342, -1, -1, 345, 346, 347, -1, -1, 350, -1, -1, 353, 354, -1, -1, 651, 358, 359, 653, 361, 362, 363, -1, -1, 366, -1, -1, 369, 655, 371, -1, -1, 374, 375, 376, 657, 378, -1, -1, 381, 382, -1, -1, 385, -1, -1, 388, 389, 659, 661, 663, 393, 394, 395, 396, 397, 398, 665, 667, 669, 402, 403, 671, 673, 406, 407, -1, -1, 675, 411, 412, 413, 677, 679, 416, 417, -1, -1, 681, 421, 422, 423, -1, -1, 683, 427, 685, 429, -1, -1, 432, 433, 434, 435, 687, 689, 438, 439, -1, -1, 442, -1, -1, 445, 446, 691, 448, -1, -1, 451, 693, 695, 454, 455, 697, 699, 458, 701, 460, 703, 462, -1, -1, 465, 466, 467, 705, 707, 470, 471, 472, 473, -1, -1, 476, -1, -1, 479, 709, 711, 482, 713, 484, 715, 717, 487, 488, 719, 490, 491, 492, -1, -1, 721, 723, 497, 725, 499, 727, 501, 502, -1, -1, 729, -1, -1, -1, -1, 731, 733, 735, 737, -1, -1, 739, 741, -1, -1, -1, -1, 743, 745, -1, -1, 747, 749, -1, -1, -1, -1, 751, 753, 755, 757, 759, 761, -1, -1, 763, 765, 767, 769, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 771, 773, -1, -1, 775, 777, 779, 781, -1, -1, -1, -1, -1, -1, 783, 785, 787, 789, 791, 793, 795, 797, 799, 801, 803, 805, 807, 809, 811, 813, 815, 817, -1, -1, 819, 821, 823, 825, -1, -1, -1, -1, -1, -1, 827, 829, 831, 833, 835, 837, 839, 841, -1, -1, -1, -1, 843, 845, -1, -1, 847, 849, -1, -1, -1, -1, 851, 853, -1, -1, 855, 857, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 859, 861, -1, -1, -1, -1, -1, -1, 863, 865, -1, -1, -1, -1, 867, 869, -1, -1, -1, -1, -1, -1, -1, -1, 871, 873, -1, -1, -1, -1, 875, 877, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 879, 881, 883, 885, 887, 889, -1, -1, 891, 893, 895, 897, -1, -1, -1, -1, 899, 901, -1, -1, -1, -1, 903, 905, -1, -1, 907, 909, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 951, 953, 955, 957, 959, 961, 963, 965, -1, -1, -1, -1, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, 1007, 1009, 1011, 1013, -1, -1, -1, -1, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, 7, 8, 9, -1, -1, 491, 13, 493, 495, 16, 17, 18, -1, -1, 497, 22, 499, 24, -1, -1, 27, 28, 29, 501, 31, -1, -1, 34, 503, 505, 37, 38, 507, 509, 511, 42, 43, 44, 45, 46, -1, -1, 513, 515, 51, 517, 53, 54, -1, -1, 519, 58, 59, 60, 61, -1, -1, 521, 65, 66, -1, -1, 523, 70, 71, 72, -1, -1, 525, 527, 77, 78, 79, 529, 81, 531, 83, 84, -1, -1, 87, -1, -1, 90, 91, 92, 93, -1, -1, 533, 535, 98, 537, 100, 539, 541, 103, 104, 105, 106, 543, 545, 547, 110, 111, 112, -1, -1, 549, 116, 117, -1, -1, 120, -1, -1, 123, 551, 125, 553, 127, 555, 129, -1, -1, 132, 133, 134, 135, 136, 137, 557, 139, -1, -1, 142, 559, 144, -1, -1, 147, 148, 149, -1, -1, 152, -1, -1, 155, 561, 563, 158, 159, 565, 161, 567, 569, 164, 165, 166, -1, -1, 169, -1, -1, 172, 571, 174, -1, -1, 177, 178, 573, 180, 575, 182, 183, -1, -1, 577, 187, 579, 189, 190, 581, 192, -1, -1, 195, 196, -1, -1, 583, 200, 201, 202, 203, 204, 585, 587, 589, 208, 591, 210, 211, -1, -1, 214, -1, -1, 593, 218, 595, 220, 221, 222, 223, -1, -1, 226, -1, -1, 229, 230, -1, -1, 597, 599, 235, 236, 237, 238, 239, 240, 241, 601, 243, -1, -1, 246, 603, 248, -1, -1, 251, 605, 253, 607, 255, -1, -1, 258, 259, 260, 261, -1, -1, 609, 265, 611, 267, -1, -1, 270, 271, 613, 615, 274, 617, 276, -1, -1, 279, 280, 281, 619, 283, 621, 623, 286, 287, 288, -1, -1, 625, 292, 627, 294, -1, -1, 297, 298, 299, 629, 301, -1, -1, 631, 305, 306, 633, 308, -1, -1, 311, 635, 313, -1, -1, 316, 637, 318, 319, 320, 321, 639, 323, -1, -1, 641, 327, 328, 329, -1, -1, 332, -1, -1, 335, 643, 337, -1, -1, 340, 341, 342, 343, -1, -1, 346, -1, -1, 349, 350, -1, -1, 645, 354, 355, 647, 357, -1, -1, 360, 361, -1, -1, 364, -1, -1, 367, 368, 369, 649, 371, 372, 373, 651, 375, -1, -1, 378, 379, -1, -1, 653, 383, 384, 385, -1, -1, 655, 389, 390, -1, -1, 393, -1, -1, 396, 397, 398, 399, 400, -1, -1, 657, 404, 405, -1, -1, 659, 409, 661, 411, 412, -1, -1, 415, -1, -1, 418, 419, 420, 663, 422, -1, -1, 665, 667, 427, 428, 429, 430, 431, 669, 671, 434, 673, 675, 437, 677, 679, 440, 441, 442, 443, -1, -1, 446, -1, -1, 449, 450, -1, -1, 453, -1, -1, 456, 457, 681, 459, -1, -1, 462, 463, -1, -1, 466, -1, -1, 469, 470, 471, 472, 473, -1, -1, 683, 477, 685, 687, 689, 481, 482, 483, 691, 485, -1, -1, 488, 693, 695, 697, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 699, 701, -1, -1, 703, 705, 707, 709, -1, -1, -1, -1, -1, -1, -1, -1, 711, 713, 715, 717, 719, 721, -1, -1, 723, 725, 727, 729, -1, -1, -1, -1, -1, -1, -1, -1, 731, 733, -1, -1, 735, 737, 739, 741, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 743, 745, -1, -1, -1, -1, -1, -1, 747, 749, 751, 753, -1, -1, 755, 757, -1, -1, -1, -1, -1, -1, -1, -1, 759, 761, 763, 765, 767, 769, 771, 773, -1, -1, 775, 777, -1, -1, -1, -1, 779, 781, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 783, 785, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 787, 789, -1, -1, -1, -1, 791, 793, -1, -1, 795, 797, -1, -1, -1, -1, -1, -1, 799, 801, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 803, 805, -1, -1, 807, 809, 811, 813, -1, -1, -1, -1, -1, -1, -1, -1, 815, 817, 819, 821, -1, -1, -1, -1, -1, -1, -1, -1, 823, 825, -1, -1, -1, -1, -1, -1, 827, 829, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 831, 833, 835, 837, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 839, 841, 843, 845, -1, -1, -1, -1, -1, -1, -1, -1, 847, 849, 851, 853, -1, -1, -1, -1, 855, 857, 859, 861, -1, -1, -1, -1, -1, -1, -1, -1, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 887, 889, 891, 893, -1, -1, -1, -1, 895, 897, 899, 901, -1, -1, -1, -1, -1, -1, -1, -1, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, 935, 937, 939, 941, 943, 945, 947, 949, 951, 953, 955, 957, -1, -1, -1, -1, -1, -1, -1, -1, 959, 961, 963, 965, 967, 969, 971, 973, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, 7, 479, 9, 10, -1, -1, 13, -1, -1, 16, 481, 483, 19, 20, 21, 485, 23, -1, -1, 26, 487, 28, -1, -1, 31, 489, 33, 491, 493, 36, 37, 38, 39, 40, -1, -1, 43, -1, -1, 495, 47, 48, 497, 50, -1, -1, 53, 499, 55, -1, -1, 58, 59, 60, 61, -1, -1, 501, 65, 66, -1, -1, 503, 70, 71, 72, -1, -1, 75, -1, -1, 505, 79, 80, 81, 507, 509, 84, 85, 86, 87, -1, -1, 511, 91, 92, -1, -1, 95, -1, -1, 98, 99, 100, -1, -1, 513, 104, 105, -1, -1, 108, -1, -1, 111, 515, 113, 114, 115, 116, -1, -1, 119, -1, -1, 122, 123, -1, -1, 126, -1, -1, 129, 130, 131, -1, -1, 134, -1, -1, 137, 138, -1, -1, 141, -1, -1, 144, 145, 146, 147, 517, 149, 519, 151, 521, 153, -1, -1, 156, 157, 158, 159, -1, -1, 523, 163, 525, 527, 529, 167, 168, 169, 170, 171, -1, -1, 531, 533, 176, 535, 178, 537, 180, -1, -1, 183, 184, 185, 539, 187, -1, -1, 541, 543, 192, 193, 194, 545, 196, 547, 198, 199, -1, -1, 202, -1, -1, 205, 549, 207, 208, 209, -1, -1, 212, -1, -1, 215, 551, 217, -1, -1, 220, 221, 222, 553, 224, 555, 557, 227, 228, 229, -1, -1, 559, 561, 234, 563, 236, 237, 565, 567, 569, 241, 242, 243, 244, 245, 246, 247, 248, -1, -1, 251, -1, -1, 571, 255, 256, 573, 258, -1, -1, 575, 262, 263, 264, 577, 266, -1, -1, 579, 270, 271, 581, 273, -1, -1, 276, 583, 278, -1, -1, 281, 585, 283, 284, 587, 589, 287, 288, 289, -1, -1, 591, 293, 294, -1, -1, 593, 298, 299, 300, 301, 302, 303, -1, -1, 595, 597, 308, 309, 599, 601, 312, 313, -1, -1, 316, -1, -1, 319, 320, 603, 322, 605, 607, 325, 609, 327, 328, -1, -1, 331, -1, -1, 334, 335, 336, 337, 338, -1, -1, 341, -1, -1, 344, 611, 346, -1, -1, 349, 350, 351, -1, -1, 613, 355, 615, 617, 358, 359, 619, 621, 623, 363, 364, 365, 625, 367, 368, 369, 627, 371, -1, -1, 629, 375, 631, 377, 633, 635, 380, 381, 382, 383, 637, 639, 386, 387, -1, -1, 390, -1, -1, 393, 394, 395, -1, -1, 398, -1, -1, 401, 402, -1, -1, 405, -1, -1, 408, 641, 410, 411, 412, -1, -1, 415, -1, -1, 418, 419, -1, -1, 422, -1, -1, 425, 426, 643, 428, 429, 430, 431, -1, -1, 434, -1, -1, 437, 438, -1, -1, 441, -1, -1, 444, 645, 446, 647, 448, -1, -1, 451, 452, 453, 454, 649, 651, 653, 655, 459, 460, 461, 462, -1, -1, 465, -1, -1, 657, 469, 470, 471, -1, -1, 659, 475, 661, 477, -1, -1, 663, 665, 667, 669, 671, 673, -1, -1, -1, -1, 675, 677, -1, -1, -1, -1, 679, 681, -1, -1, -1, -1, -1, -1, -1, -1, 683, 685, 687, 689, 691, 693, -1, -1, -1, -1, 695, 697, 699, 701, 703, 705, -1, -1, -1, -1, -1, -1, -1, -1, 707, 709, -1, -1, 711, 713, 715, 717, -1, -1, -1, -1, 719, 721, 723, 725, 727, 729, 731, 733, 735, 737, -1, -1, 739, 741, -1, -1, -1, -1, -1, -1, 743, 745, 747, 749, -1, -1, -1, -1, 751, 753, 755, 757, -1, -1, 759, 761, -1, -1, 763, 765, -1, -1, -1, -1, 767, 769, 771, 773, 775, 777, -1, -1, -1, -1, -1, -1, 779, 781, -1, -1, -1, -1, 783, 785, -1, -1, -1, -1, 787, 789, -1, -1, -1, -1, -1, -1, -1, -1, 791, 793, 795, 797, 799, 801, 803, 805, -1, -1, 807, 809, 811, 813, -1, -1, -1, -1, -1, -1, -1, -1, 815, 817, 819, 821, 823, 825, -1, -1, -1, -1, -1, -1, 827, 829, 831, 833, 835, 837, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 839, 841, 843, 845, 847, 849, 851, 853, 855, 857, 859, 861, 863, 865, 867, 869, -1, -1, -1, -1, 871, 873, 875, 877, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 879, 881, 883, 885, 887, 889, 891, 893, -1, -1, -1, -1, 895, 897, 899, 901, -1, -1, -1, -1, -1, -1, -1, -1, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, 943, 945, 947, 949, -1, -1, -1, -1, -1, -1, -1, -1, 951, 953, 955, 957, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 959, 961, 963, 965, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((230, 137, 86, 33, 18, 11, 10, 9, 506, 508, 510, 13, 512, 15, 514, 17, -1, -1, 28, 21, 516, 25, 24, -1, -1, 27, -1, -1, 32, 31, 518, 520, 522, 57, 48, 41, 38, 524, 40, -1, -1, 45, 44, -1, -1, 47, -1, -1, 56, 53, 52, -1, -1, 55, -1, -1, 526, 71, 66, 63, 62, -1, -1, 65, -1, -1, 68, 528, 70, -1, -1, 79, 76, 75, -1, -1, 78, -1, -1, 83, 82, -1, -1, 85, -1, -1, 106, 97, 96, 95, 94, 93, -1, -1, 530, 532, 534, 99, 536, 105, 102, 538, 104, -1, -1, 540, 124, 113, 110, 542, 112, 544, 546, 119, 118, 117, -1, -1, 548, 123, 122, -1, -1, 550, 130, 129, 128, 552, 554, 556, 136, 135, 134, -1, -1, 558, 560, 189, 164, 159, 148, 143, 562, 145, 564, 147, -1, -1, 154, 151, 566, 153, -1, -1, 156, 568, 158, -1, -1, 163, 162, 570, 572, 574, 176, 175, 174, 171, 170, -1, -1, 173, -1, -1, 576, 578, 186, 185, 182, 181, -1, -1, 184, -1, -1, 580, 188, 582, 584, 211, 200, 199, 194, 586, 196, 588, 198, -1, -1, 590, 202, 592, 206, 205, 594, 596, 208, 598, 210, -1, -1, 217, 216, 215, 600, 602, 604, 223, 220, 606, 222, 608, 610, 225, 612, 229, 228, -1, -1, 614, 392, 315, 266, 247, 240, 237, 616, 239, 618, 620, 242, 622, 244, 624, 246, -1, -1, 255, 250, 626, 252, 628, 254, -1, -1, 261, 258, 630, 260, -1, -1, 265, 264, -1, -1, 632, 294, 281, 276, 273, 272, -1, -1, 275, -1, -1, 280, 279, -1, -1, 634, 287, 286, 285, -1, -1, 636, 291, 290, -1, -1, 293, -1, -1, 302, 301, 298, 638, 300, -1, -1, 640, 308, 305, 642, 307, -1, -1, 312, 311, -1, -1, 314, -1, -1, 357, 330, 329, 324, 321, 644, 323, -1, -1, 326, 646, 328, -1, -1, 648, 344, 337, 336, 335, -1, -1, 650, 341, 340, -1, -1, 343, -1, -1, 352, 349, 348, -1, -1, 351, -1, -1, 356, 355, -1, -1, 652, 373, 360, 654, 368, 365, 364, -1, -1, 367, -1, -1, 370, 656, 372, -1, -1, 387, 380, 377, 658, 379, -1, -1, 384, 383, -1, -1, 386, -1, -1, 391, 390, 660, 662, 664, 464, 431, 410, 401, 400, 399, 666, 668, 670, 405, 404, 672, 674, 409, 408, -1, -1, 676, 420, 415, 414, 678, 680, 419, 418, -1, -1, 682, 426, 425, 424, -1, -1, 684, 428, 686, 430, -1, -1, 453, 444, 437, 436, 688, 690, 441, 440, -1, -1, 443, -1, -1, 450, 447, 692, 449, -1, -1, 452, 694, 696, 457, 456, 698, 700, 459, 702, 461, 704, 463, -1, -1, 486, 469, 468, 706, 708, 481, 478, 475, 474, -1, -1, 477, -1, -1, 480, 710, 712, 483, 714, 485, 716, 718, 496, 489, 720, 495, 494, 493, -1, -1, 722, 724, 498, 726, 500, 728, 504, 503, -1, -1, 730, -1, -1, -1, -1, 732, 734, 736, 738, -1, -1, 740, 742, -1, -1, -1, -1, 744, 746, -1, -1, 748, 750, -1, -1, -1, -1, 752, 754, 756, 758, 760, 762, -1, -1, 764, 766, 768, 770, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 772, 774, -1, -1, 776, 778, 780, 782, -1, -1, -1, -1, -1, -1, 784, 786, 788, 790, 792, 794, 796, 798, 800, 802, 804, 806, 808, 810, 812, 814, 816, 818, -1, -1, 820, 822, 824, 826, -1, -1, -1, -1, -1, -1, 828, 830, 832, 834, 836, 838, 840, 842, -1, -1, -1, -1, 844, 846, -1, -1, 848, 850, -1, -1, -1, -1, 852, 854, -1, -1, 856, 858, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 860, 862, -1, -1, -1, -1, -1, -1, 864, 866, -1, -1, -1, -1, 868, 870, -1, -1, -1, -1, -1, -1, -1, -1, 872, 874, -1, -1, -1, -1, 876, 878, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 880, 882, 884, 886, 888, 890, -1, -1, 892, 894, 896, 898, -1, -1, -1, -1, 900, 902, -1, -1, -1, -1, 904, 906, -1, -1, 908, 910, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 952, 954, 956, 958, 960, 962, 964, 966, -1, -1, -1, -1, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, 1008, 1010, 1012, 1014, -1, -1, -1, -1, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (234, 131, 76, 41, 26, 15, 12, 11, 10, -1, -1, 492, 14, 494, 496, 21, 20, 19, -1, -1, 498, 23, 500, 25, -1, -1, 36, 33, 30, 502, 32, -1, -1, 35, 504, 506, 40, 39, 508, 510, 512, 57, 50, 49, 48, 47, -1, -1, 514, 516, 52, 518, 56, 55, -1, -1, 520, 69, 64, 63, 62, -1, -1, 522, 68, 67, -1, -1, 524, 75, 74, 73, -1, -1, 526, 528, 102, 89, 80, 530, 82, 532, 86, 85, -1, -1, 88, -1, -1, 97, 96, 95, 94, -1, -1, 534, 536, 99, 538, 101, 540, 542, 122, 109, 108, 107, 544, 546, 548, 115, 114, 113, -1, -1, 550, 119, 118, -1, -1, 121, -1, -1, 124, 552, 126, 554, 128, 556, 130, -1, -1, 199, 176, 157, 146, 141, 138, 558, 140, -1, -1, 143, 560, 145, -1, -1, 154, 151, 150, -1, -1, 153, -1, -1, 156, 562, 564, 163, 160, 566, 162, 568, 570, 171, 168, 167, -1, -1, 170, -1, -1, 173, 572, 175, -1, -1, 186, 179, 574, 181, 576, 185, 184, -1, -1, 578, 188, 580, 194, 191, 582, 193, -1, -1, 198, 197, -1, -1, 584, 217, 216, 207, 206, 205, 586, 588, 590, 209, 592, 213, 212, -1, -1, 215, -1, -1, 594, 219, 596, 233, 228, 225, 224, -1, -1, 227, -1, -1, 232, 231, -1, -1, 598, 600, 366, 315, 278, 257, 250, 245, 242, 602, 244, -1, -1, 247, 604, 249, -1, -1, 252, 606, 254, 608, 256, -1, -1, 269, 264, 263, 262, -1, -1, 610, 266, 612, 268, -1, -1, 273, 272, 614, 616, 275, 618, 277, -1, -1, 296, 285, 282, 620, 284, 622, 624, 291, 290, 289, -1, -1, 626, 293, 628, 295, -1, -1, 304, 303, 300, 630, 302, -1, -1, 632, 310, 307, 634, 309, -1, -1, 312, 636, 314, -1, -1, 317, 638, 339, 326, 325, 322, 640, 324, -1, -1, 642, 334, 331, 330, -1, -1, 333, -1, -1, 336, 644, 338, -1, -1, 353, 348, 345, 344, -1, -1, 347, -1, -1, 352, 351, -1, -1, 646, 359, 356, 648, 358, -1, -1, 363, 362, -1, -1, 365, -1, -1, 426, 395, 370, 650, 382, 377, 374, 652, 376, -1, -1, 381, 380, -1, -1, 654, 388, 387, 386, -1, -1, 656, 392, 391, -1, -1, 394, -1, -1, 417, 408, 403, 402, 401, -1, -1, 658, 407, 406, -1, -1, 660, 410, 662, 414, 413, -1, -1, 416, -1, -1, 425, 424, 421, 664, 423, -1, -1, 666, 668, 468, 439, 436, 433, 432, 670, 672, 435, 674, 676, 438, 678, 680, 455, 448, 445, 444, -1, -1, 447, -1, -1, 452, 451, -1, -1, 454, -1, -1, 461, 458, 682, 460, -1, -1, 465, 464, -1, -1, 467, -1, -1, 480, 479, 476, 475, 474, -1, -1, 684, 478, 686, 688, 690, 490, 487, 484, 692, 486, -1, -1, 489, 694, 696, 698, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 700, 702, -1, -1, 704, 706, 708, 710, -1, -1, -1, -1, -1, -1, -1, -1, 712, 714, 716, 718, 720, 722, -1, -1, 724, 726, 728, 730, -1, -1, -1, -1, -1, -1, -1, -1, 732, 734, -1, -1, 736, 738, 740, 742, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 744, 746, -1, -1, -1, -1, -1, -1, 748, 750, 752, 754, -1, -1, 756, 758, -1, -1, -1, -1, -1, -1, -1, -1, 760, 762, 764, 766, 768, 770, 772, 774, -1, -1, 776, 778, -1, -1, -1, -1, 780, 782, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 784, 786, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 788, 790, -1, -1, -1, -1, 792, 794, -1, -1, 796, 798, -1, -1, -1, -1, -1, -1, 800, 802, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 804, 806, -1, -1, 808, 810, 812, 814, -1, -1, -1, -1, -1, -1, -1, -1, 816, 818, 820, 822, -1, -1, -1, -1, -1, -1, -1, -1, 824, 826, -1, -1, -1, -1, -1, -1, 828, 830, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 832, 834, 836, 838, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 840, 842, 844, 846, -1, -1, -1, -1, -1, -1, -1, -1, 848, 850, 852, 854, -1, -1, -1, -1, 856, 858, 860, 862, -1, -1, -1, -1, -1, -1, -1, -1, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 888, 890, 892, 894, -1, -1, -1, -1, 896, 898, 900, 902, -1, -1, -1, -1, -1, -1, -1, -1, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, 936, 938, 940, 942, 944, 946, 948, 950, 952, 954, 956, 958, -1, -1, -1, -1, -1, -1, -1, -1, 960, 962, 964, 966, 968, 970, 972, 974, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (240, 143, 78, 35, 18, 15, 8, 480, 12, 11, -1, -1, 14, -1, -1, 17, 482, 484, 30, 25, 22, 486, 24, -1, -1, 27, 488, 29, -1, -1, 32, 490, 34, 492, 494, 57, 46, 45, 42, 41, -1, -1, 44, -1, -1, 496, 52, 49, 498, 51, -1, -1, 54, 500, 56, -1, -1, 69, 64, 63, 62, -1, -1, 502, 68, 67, -1, -1, 504, 77, 74, 73, -1, -1, 76, -1, -1, 506, 110, 83, 82, 508, 510, 97, 90, 89, 88, -1, -1, 512, 94, 93, -1, -1, 96, -1, -1, 103, 102, 101, -1, -1, 514, 107, 106, -1, -1, 109, -1, -1, 112, 516, 128, 121, 118, 117, -1, -1, 120, -1, -1, 125, 124, -1, -1, 127, -1, -1, 136, 133, 132, -1, -1, 135, -1, -1, 140, 139, -1, -1, 142, -1, -1, 191, 166, 155, 148, 518, 150, 520, 152, 522, 154, -1, -1, 165, 162, 161, 160, -1, -1, 524, 164, 526, 528, 530, 182, 175, 174, 173, 172, -1, -1, 532, 534, 177, 536, 179, 538, 181, -1, -1, 190, 189, 186, 540, 188, -1, -1, 542, 544, 219, 204, 195, 546, 197, 548, 201, 200, -1, -1, 203, -1, -1, 206, 550, 214, 211, 210, -1, -1, 213, -1, -1, 216, 552, 218, -1, -1, 233, 226, 223, 554, 225, 556, 558, 232, 231, 230, -1, -1, 560, 562, 235, 564, 239, 238, 566, 568, 570, 362, 297, 280, 261, 254, 253, 250, 249, -1, -1, 252, -1, -1, 572, 260, 257, 574, 259, -1, -1, 576, 269, 268, 265, 578, 267, -1, -1, 580, 275, 272, 582, 274, -1, -1, 277, 584, 279, -1, -1, 282, 586, 286, 285, 588, 590, 292, 291, 290, -1, -1, 592, 296, 295, -1, -1, 594, 333, 318, 307, 306, 305, 304, -1, -1, 596, 598, 311, 310, 600, 602, 315, 314, -1, -1, 317, -1, -1, 324, 321, 604, 323, 606, 608, 326, 610, 330, 329, -1, -1, 332, -1, -1, 357, 348, 343, 340, 339, -1, -1, 342, -1, -1, 345, 612, 347, -1, -1, 354, 353, 352, -1, -1, 614, 356, 616, 618, 361, 360, 620, 622, 624, 424, 379, 366, 626, 374, 373, 370, 628, 372, -1, -1, 630, 376, 632, 378, 634, 636, 407, 392, 385, 384, 638, 640, 389, 388, -1, -1, 391, -1, -1, 400, 397, 396, -1, -1, 399, -1, -1, 404, 403, -1, -1, 406, -1, -1, 409, 642, 417, 414, 413, -1, -1, 416, -1, -1, 421, 420, -1, -1, 423, -1, -1, 450, 427, 644, 443, 436, 433, 432, -1, -1, 435, -1, -1, 440, 439, -1, -1, 442, -1, -1, 445, 646, 447, 648, 449, -1, -1, 458, 457, 456, 455, 650, 652, 654, 656, 468, 467, 464, 463, -1, -1, 466, -1, -1, 658, 474, 473, 472, -1, -1, 660, 476, 662, 478, -1, -1, 664, 666, 668, 670, 672, 674, -1, -1, -1, -1, 676, 678, -1, -1, -1, -1, 680, 682, -1, -1, -1, -1, -1, -1, -1, -1, 684, 686, 688, 690, 692, 694, -1, -1, -1, -1, 696, 698, 700, 702, 704, 706, -1, -1, -1, -1, -1, -1, -1, -1, 708, 710, -1, -1, 712, 714, 716, 718, -1, -1, -1, -1, 720, 722, 724, 726, 728, 730, 732, 734, 736, 738, -1, -1, 740, 742, -1, -1, -1, -1, -1, -1, 744, 746, 748, 750, -1, -1, -1, -1, 752, 754, 756, 758, -1, -1, 760, 762, -1, -1, 764, 766, -1, -1, -1, -1, 768, 770, 772, 774, 776, 778, -1, -1, -1, -1, -1, -1, 780, 782, -1, -1, -1, -1, 784, 786, -1, -1, -1, -1, 788, 790, -1, -1, -1, -1, -1, -1, -1, -1, 792, 794, 796, 798, 800, 802, 804, 806, -1, -1, 808, 810, 812, 814, -1, -1, -1, -1, -1, -1, -1, -1, 816, 818, 820, 822, 824, 826, -1, -1, -1, -1, -1, -1, 828, 830, 832, 834, 836, 838, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 840, 842, 844, 846, 848, 850, 852, 854, 856, 858, 860, 862, 864, 866, 868, 870, -1, -1, -1, -1, 872, 874, 876, 878, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 880, 882, 884, 886, 888, 890, 892, 894, -1, -1, -1, -1, 896, 898, 900, 902, -1, -1, -1, -1, -1, -1, -1, -1, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, 944, 946, 948, 950, -1, -1, -1, -1, -1, -1, -1, -1, 952, 954, 956, 958, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 960, 962, 964, 966, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 1, 2, 3, 4, 5, 6, 7, 7, 6, 5, 11, 11, 13, 13, 15, 15, 4, 18, 19, 19, 21, 22, 22, 21, 25, 25, 18, 28, 29, 29, 28, 3, 33, 34, 35, 36, 36, 38, 38, 35, 41, 42, 42, 41, 45, 45, 34, 48, 49, 50, 50, 49, 53, 53, 48, 33, 57, 58, 59, 60, 60, 59, 63, 63, 58, 66, 66, 68, 68, 57, 71, 72, 73, 73, 72, 76, 76, 71, 79, 80, 80, 79, 83, 83, 2, 86, 87, 88, 89, 90, 91, 91, 90, 89, 88, 87, 97, 97, 99, 100, 100, 102, 102, 99, 86, 106, 107, 108, 108, 110, 110, 107, 113, 114, 115, 115, 114, 113, 119, 120, 120, 119, 106, 124, 125, 126, 126, 125, 124, 130, 131, 132, 132, 131, 130, 1, 137, 138, 139, 140, 141, 141, 143, 143, 145, 145, 140, 148, 149, 149, 151, 151, 148, 154, 154, 156, 156, 139, 159, 160, 160, 159, 138, 164, 165, 166, 167, 168, 168, 167, 171, 171, 166, 165, 164, 176, 177, 178, 179, 179, 178, 182, 182, 177, 176, 186, 186, 137, 189, 190, 191, 192, 192, 194, 194, 196, 196, 191, 190, 200, 200, 202, 203, 203, 202, 206, 206, 208, 208, 189, 211, 212, 213, 213, 212, 211, 217, 218, 218, 220, 220, 217, 223, 223, 225, 226, 226, 225, 0, 230, 231, 232, 233, 234, 235, 235, 237, 237, 234, 240, 240, 242, 242, 244, 244, 233, 247, 248, 248, 250, 250, 252, 252, 247, 255, 256, 256, 258, 258, 255, 261, 262, 262, 261, 232, 266, 267, 268, 269, 270, 270, 269, 273, 273, 268, 276, 277, 277, 276, 267, 281, 282, 283, 283, 282, 281, 287, 288, 288, 287, 291, 291, 266, 294, 295, 296, 296, 298, 298, 295, 294, 302, 303, 303, 305, 305, 302, 308, 309, 309, 308, 312, 312, 231, 315, 316, 317, 318, 319, 319, 321, 321, 318, 324, 324, 326, 326, 317, 316, 330, 331, 332, 333, 333, 332, 331, 337, 338, 338, 337, 341, 341, 330, 344, 345, 346, 346, 345, 349, 349, 344, 352, 353, 353, 352, 315, 357, 358, 358, 360, 361, 362, 362, 361, 365, 365, 360, 368, 368, 370, 370, 357, 373, 374, 375, 375, 377, 377, 374, 380, 381, 381, 380, 384, 384, 373, 387, 388, 388, 387, 230, 392, 393, 394, 395, 396, 397, 397, 396, 395, 401, 402, 402, 401, 405, 406, 406, 405, 394, 410, 411, 412, 412, 411, 415, 416, 416, 415, 410, 420, 421, 422, 422, 421, 420, 426, 426, 428, 428, 393, 431, 432, 433, 434, 434, 433, 437, 438, 438, 437, 441, 441, 432, 444, 445, 445, 447, 447, 444, 450, 450, 431, 453, 454, 454, 453, 457, 457, 459, 459, 461, 461, 392, 464, 465, 466, 466, 465, 469, 470, 471, 472, 472, 471, 475, 475, 470, 478, 478, 469, 481, 481, 483, 483, 464, 486, 487, 487, 489, 490, 491, 491, 490, 489, 486, 496, 496, 498, 498, 500, 501, 501, 500, 8, 8, 9, 9, 10, 10, 12, 12, 14, 14, 20, 20, 30, 30, 31, 31, 32, 32, 37, 37, 56, 56, 67, 67, 94, 94, 95, 95, 96, 96, 98, 98, 101, 101, 105, 105, 109, 109, 111, 111, 112, 112, 118, 118, 123, 123, 127, 127, 128, 128, 129, 129, 135, 135, 136, 136, 142, 142, 144, 144, 150, 150, 155, 155, 161, 161, 162, 162, 163, 163, 174, 174, 175, 175, 185, 185, 187, 187, 188, 188, 193, 193, 195, 195, 199, 199, 201, 201, 204, 204, 205, 205, 207, 207, 214, 214, 215, 215, 216, 216, 219, 219, 221, 221, 222, 222, 224, 224, 229, 229, 236, 236, 238, 238, 239, 239, 241, 241, 243, 243, 249, 249, 251, 251, 257, 257, 265, 265, 280, 280, 286, 286, 297, 297, 301, 301, 304, 304, 320, 320, 325, 325, 329, 329, 336, 336, 356, 356, 359, 359, 369, 369, 376, 376, 389, 389, 390, 390, 391, 391, 398, 398, 399, 399, 400, 400, 403, 403, 404, 404, 409, 409, 413, 413, 414, 414, 419, 419, 425, 425, 427, 427, 435, 435, 436, 436, 446, 446, 451, 451, 452, 452, 455, 455, 456, 456, 458, 458, 460, 460, 467, 467, 468, 468, 479, 479, 480, 480, 482, 482, 484, 484, 485, 485, 488, 488, 494, 494, 495, 495, 497, 497, 499, 499, 504, 504, 509, 509, 510, 510, 511, 511, 512, 512, 515, 515, 516, 516, 521, 521, 522, 522, 525, 525, 526, 526, 531, 531, 532, 532, 533, 533, 534, 534, 535, 535, 536, 536, 539, 539, 540, 540, 541, 541, 542, 542, 555, 555, 556, 556, 559, 559, 560, 560, 561, 561, 562, 562, 569, 569, 570, 570, 571, 571, 572, 572, 573, 573, 574, 574, 575, 575, 576, 576, 577, 577, 578, 578, 579, 579, 580, 580, 581, 581, 582, 582, 583, 583, 584, 584, 585, 585, 586, 586, 589, 589, 590, 590, 591, 591, 592, 592, 599, 599, 600, 600, 601, 601, 602, 602, 603, 603, 604, 604, 605, 605, 606, 606, 611, 611, 612, 612, 615, 615, 616, 616, 621, 621, 622, 622, 625, 625, 626, 626, 639, 639, 640, 640, 647, 647, 648, 648, 653, 653, 654, 654, 663, 663, 664, 664, 669, 669, 670, 670, 697, 697, 698, 698, 699, 699, 700, 700, 701, 701, 702, 702, 705, 705, 706, 706, 707, 707, 708, 708, 713, 713, 714, 714, 719, 719, 720, 720, 723, 723, 724, 724, 725, 725, 726, 726, 727, 727, 728, 728, 755, 755, 756, 756, 757, 757, 758, 758, 759, 759, 760, 760, 761, 761, 762, 762, 791, 791, 792, 792, 793, 793, 794, 794, 799, 799, 800, 800, 801, 801, 802, 802, 819, 819, 820, 820, 821, 821, 822, 822, 823, 823, 824, 824, 825, 825, 826, 826, 835, 835, 836, 836, 837, 837, 838, 838, 863, 863, 864, 864, 865, 865, 866, 866, 867, 867, 868, 868, 869, 869, 870, 870, 891, 891, 892, 892, 893, 893, 894, 894, 895, 895, 896, 896, 897, 897, 898, 898, 903, 903, 904, 904, 905, 905, 906, 906, 911, 911, 912, 912, 913, 913, 914, 914),
                (-1, 0, 1, 2, 3, 4, 5, 6, 7, 8, 8, 7, 6, 12, 12, 5, 15, 16, 17, 17, 16, 15, 21, 21, 23, 23, 4, 26, 27, 28, 28, 30, 30, 27, 33, 33, 26, 36, 37, 37, 36, 3, 41, 42, 43, 44, 45, 45, 44, 43, 42, 50, 50, 52, 53, 53, 52, 41, 57, 58, 59, 60, 60, 59, 58, 64, 65, 65, 64, 57, 69, 70, 71, 71, 70, 69, 2, 76, 77, 78, 78, 80, 80, 82, 83, 83, 82, 86, 86, 77, 89, 90, 91, 92, 92, 91, 90, 89, 97, 97, 99, 99, 76, 102, 103, 104, 105, 105, 104, 103, 109, 110, 111, 111, 110, 109, 115, 116, 116, 115, 119, 119, 102, 122, 122, 124, 124, 126, 126, 128, 128, 1, 131, 132, 133, 134, 135, 136, 136, 138, 138, 135, 141, 141, 143, 143, 134, 146, 147, 148, 148, 147, 151, 151, 146, 154, 154, 133, 157, 158, 158, 160, 160, 157, 163, 164, 165, 165, 164, 168, 168, 163, 171, 171, 173, 173, 132, 176, 177, 177, 179, 179, 181, 182, 182, 181, 176, 186, 186, 188, 189, 189, 191, 191, 188, 194, 195, 195, 194, 131, 199, 200, 201, 202, 203, 203, 202, 201, 207, 207, 209, 210, 210, 209, 213, 213, 200, 199, 217, 217, 219, 220, 221, 222, 222, 221, 225, 225, 220, 228, 229, 229, 228, 219, 0, 234, 235, 236, 237, 238, 239, 240, 240, 242, 242, 239, 245, 245, 247, 247, 238, 250, 250, 252, 252, 254, 254, 237, 257, 258, 259, 260, 260, 259, 258, 264, 264, 266, 266, 257, 269, 270, 270, 269, 273, 273, 275, 275, 236, 278, 279, 280, 280, 282, 282, 279, 285, 286, 287, 287, 286, 285, 291, 291, 293, 293, 278, 296, 297, 298, 298, 300, 300, 297, 296, 304, 305, 305, 307, 307, 304, 310, 310, 312, 312, 235, 315, 315, 317, 318, 319, 320, 320, 322, 322, 319, 318, 326, 327, 328, 328, 327, 331, 331, 326, 334, 334, 336, 336, 317, 339, 340, 341, 342, 342, 341, 345, 345, 340, 348, 349, 349, 348, 339, 353, 354, 354, 356, 356, 353, 359, 360, 360, 359, 363, 363, 234, 366, 367, 368, 368, 370, 371, 372, 372, 374, 374, 371, 377, 378, 378, 377, 370, 382, 383, 384, 384, 383, 382, 388, 389, 389, 388, 392, 392, 367, 395, 396, 397, 398, 399, 399, 398, 397, 403, 404, 404, 403, 396, 408, 408, 410, 411, 411, 410, 414, 414, 395, 417, 418, 419, 419, 421, 421, 418, 417, 366, 426, 427, 428, 429, 430, 430, 429, 433, 433, 428, 436, 436, 427, 439, 440, 441, 442, 442, 441, 445, 445, 440, 448, 449, 449, 448, 452, 452, 439, 455, 456, 456, 458, 458, 455, 461, 462, 462, 461, 465, 465, 426, 468, 469, 470, 471, 472, 472, 471, 470, 476, 476, 469, 468, 480, 481, 482, 482, 484, 484, 481, 487, 487, 480, 11, 11, 13, 13, 14, 14, 20, 20, 22, 22, 29, 29, 34, 34, 35, 35, 38, 38, 39, 39, 40, 40, 48, 48, 49, 49, 51, 51, 56, 56, 63, 63, 68, 68, 74, 74, 75, 75, 79, 79, 81, 81, 95, 95, 96, 96, 98, 98, 100, 100, 101, 101, 106, 106, 107, 107, 108, 108, 114, 114, 123, 123, 125, 125, 127, 127, 137, 137, 142, 142, 155, 155, 156, 156, 159, 159, 161, 161, 162, 162, 172, 172, 178, 178, 180, 180, 185, 185, 187, 187, 190, 190, 198, 198, 204, 204, 205, 205, 206, 206, 208, 208, 216, 216, 218, 218, 232, 232, 233, 233, 241, 241, 246, 246, 251, 251, 253, 253, 263, 263, 265, 265, 271, 271, 272, 272, 274, 274, 281, 281, 283, 283, 284, 284, 290, 290, 292, 292, 299, 299, 303, 303, 306, 306, 311, 311, 316, 316, 321, 321, 325, 325, 335, 335, 352, 352, 355, 355, 369, 369, 373, 373, 381, 381, 387, 387, 402, 402, 407, 407, 409, 409, 420, 420, 424, 424, 425, 425, 431, 431, 432, 432, 434, 434, 435, 435, 437, 437, 438, 438, 457, 457, 475, 475, 477, 477, 478, 478, 479, 479, 483, 483, 488, 488, 489, 489, 490, 490, 511, 511, 512, 512, 515, 515, 516, 516, 517, 517, 518, 518, 527, 527, 528, 528, 529, 529, 530, 530, 531, 531, 532, 532, 535, 535, 536, 536, 537, 537, 538, 538, 547, 547, 548, 548, 551, 551, 552, 552, 553, 553, 554, 554, 565, 565, 566, 566, 573, 573, 574, 574, 575, 575, 576, 576, 579, 579, 580, 580, 589, 589, 590, 590, 591, 591, 592, 592, 593, 593, 594, 594, 595, 595, 596, 596, 599, 599, 600, 600, 605, 605, 606, 606, 619, 619, 620, 620, 631, 631, 632, 632, 637, 637, 638, 638, 641, 641, 642, 642, 649, 649, 650, 650, 661, 661, 662, 662, 665, 665, 666, 666, 667, 667, 668, 668, 677, 677, 678, 678, 679, 679, 680, 680, 689, 689, 690, 690, 697, 697, 698, 698, 715, 715, 716, 716, 717, 717, 718, 718, 735, 735, 736, 736, 737, 737, 738, 738, 747, 747, 748, 748, 749, 749, 750, 750, 755, 755, 756, 756, 757, 757, 758, 758, 767, 767, 768, 768, 769, 769, 770, 770, 771, 771, 772, 772, 773, 773, 774, 774, 775, 775, 776, 776, 777, 777, 778, 778, 791, 791, 792, 792, 793, 793, 794, 794, 799, 799, 800, 800, 801, 801, 802, 802, 811, 811, 812, 812, 813, 813, 814, 814, 823, 823, 824, 824, 825, 825, 826, 826, 827, 827, 828, 828, 829, 829, 830, 830, 863, 863, 864, 864, 865, 865, 866, 866, 867, 867, 868, 868, 869, 869, 870, 870, 871, 871, 872, 872, 873, 873, 874, 874, 875, 875, 876, 876, 877, 877, 878, 878, 887, 887, 888, 888, 889, 889, 890, 890, 891, 891, 892, 892, 893, 893, 894, 894, 895, 895, 896, 896, 897, 897, 898, 898, 899, 899, 900, 900, 901, 901, 902, 902, 959, 959, 960, 960, 961, 961, 962, 962, 963, 963, 964, 964, 965, 965, 966, 966, 967, 967, 968, 968, 969, 969, 970, 970, 971, 971, 972, 972, 973, 973, 974, 974),
                (-1, 0, 1, 2, 3, 4, 5, 6, 6, 8, 9, 9, 8, 12, 12, 5, 15, 15, 4, 18, 19, 20, 20, 22, 22, 19, 25, 25, 27, 27, 18, 30, 30, 32, 32, 3, 35, 36, 37, 38, 39, 39, 38, 42, 42, 37, 36, 46, 47, 47, 49, 49, 46, 52, 52, 54, 54, 35, 57, 58, 59, 60, 60, 59, 58, 64, 65, 65, 64, 57, 69, 70, 71, 71, 70, 74, 74, 69, 2, 78, 79, 80, 80, 79, 83, 84, 85, 86, 86, 85, 84, 90, 91, 91, 90, 94, 94, 83, 97, 98, 99, 99, 98, 97, 103, 104, 104, 103, 107, 107, 78, 110, 110, 112, 113, 114, 115, 115, 114, 118, 118, 113, 121, 122, 122, 121, 125, 125, 112, 128, 129, 130, 130, 129, 133, 133, 128, 136, 137, 137, 136, 140, 140, 1, 143, 144, 145, 146, 146, 148, 148, 150, 150, 152, 152, 145, 155, 156, 157, 158, 158, 157, 156, 162, 162, 155, 144, 166, 167, 168, 169, 170, 170, 169, 168, 167, 175, 175, 177, 177, 179, 179, 166, 182, 183, 184, 184, 186, 186, 183, 182, 143, 191, 192, 193, 193, 195, 195, 197, 198, 198, 197, 201, 201, 192, 204, 204, 206, 207, 208, 208, 207, 211, 211, 206, 214, 214, 216, 216, 191, 219, 220, 221, 221, 223, 223, 220, 226, 227, 228, 228, 227, 226, 219, 233, 233, 235, 236, 236, 235, 0, 240, 241, 242, 243, 244, 245, 246, 247, 247, 246, 250, 250, 245, 244, 254, 255, 255, 257, 257, 254, 243, 261, 262, 263, 263, 265, 265, 262, 261, 269, 270, 270, 272, 272, 269, 275, 275, 277, 277, 242, 280, 280, 282, 283, 283, 282, 286, 287, 288, 288, 287, 286, 292, 293, 293, 292, 241, 297, 298, 299, 300, 301, 302, 302, 301, 300, 299, 307, 308, 308, 307, 311, 312, 312, 311, 315, 315, 298, 318, 319, 319, 321, 321, 318, 324, 324, 326, 327, 327, 326, 330, 330, 297, 333, 334, 335, 336, 337, 337, 336, 340, 340, 335, 343, 343, 345, 345, 334, 348, 349, 350, 350, 349, 348, 354, 354, 333, 357, 358, 358, 357, 240, 362, 363, 364, 364, 366, 367, 368, 368, 370, 370, 367, 366, 374, 374, 376, 376, 363, 379, 380, 381, 382, 382, 381, 385, 386, 386, 385, 389, 389, 380, 392, 393, 394, 394, 393, 397, 397, 392, 400, 401, 401, 400, 404, 404, 379, 407, 407, 409, 410, 411, 411, 410, 414, 414, 409, 417, 418, 418, 417, 421, 421, 362, 424, 425, 425, 427, 428, 429, 430, 430, 429, 433, 433, 428, 436, 437, 437, 436, 440, 440, 427, 443, 443, 445, 445, 447, 447, 424, 450, 451, 452, 453, 453, 452, 451, 450, 458, 459, 460, 461, 461, 460, 464, 464, 459, 458, 468, 469, 470, 470, 469, 468, 474, 474, 476, 476, 7, 7, 16, 16, 17, 17, 21, 21, 26, 26, 31, 31, 33, 33, 34, 34, 45, 45, 48, 48, 53, 53, 63, 63, 68, 68, 77, 77, 81, 81, 82, 82, 89, 89, 102, 102, 111, 111, 147, 147, 149, 149, 151, 151, 161, 161, 163, 163, 164, 164, 165, 165, 173, 173, 174, 174, 176, 176, 178, 178, 185, 185, 189, 189, 190, 190, 194, 194, 196, 196, 205, 205, 215, 215, 222, 222, 224, 224, 225, 225, 231, 231, 232, 232, 234, 234, 237, 237, 238, 238, 239, 239, 253, 253, 256, 256, 260, 260, 264, 264, 268, 268, 271, 271, 276, 276, 281, 281, 284, 284, 285, 285, 291, 291, 296, 296, 305, 305, 306, 306, 309, 309, 310, 310, 320, 320, 322, 322, 323, 323, 325, 325, 344, 344, 353, 353, 355, 355, 356, 356, 359, 359, 360, 360, 361, 361, 365, 365, 369, 369, 373, 373, 375, 375, 377, 377, 378, 378, 383, 383, 384, 384, 408, 408, 426, 426, 444, 444, 446, 446, 454, 454, 455, 455, 456, 456, 457, 457, 467, 467, 473, 473, 475, 475, 479, 479, 480, 480, 481, 481, 482, 482, 483, 483, 484, 484, 489, 489, 490, 490, 495, 495, 496, 496, 505, 505, 506, 506, 507, 507, 508, 508, 509, 509, 510, 510, 515, 515, 516, 516, 517, 517, 518, 518, 519, 519, 520, 520, 529, 529, 530, 530, 533, 533, 534, 534, 535, 535, 536, 536, 541, 541, 542, 542, 543, 543, 544, 544, 545, 545, 546, 546, 547, 547, 548, 548, 549, 549, 550, 550, 553, 553, 554, 554, 561, 561, 562, 562, 563, 563, 564, 564, 569, 569, 570, 570, 571, 571, 572, 572, 575, 575, 576, 576, 579, 579, 580, 580, 585, 585, 586, 586, 587, 587, 588, 588, 589, 589, 590, 590, 597, 597, 598, 598, 603, 603, 604, 604, 609, 609, 610, 610, 619, 619, 620, 620, 621, 621, 622, 622, 623, 623, 624, 624, 625, 625, 626, 626, 629, 629, 630, 630, 631, 631, 632, 632, 641, 641, 642, 642, 643, 643, 644, 644, 645, 645, 646, 646, 653, 653, 654, 654, 655, 655, 656, 656, 657, 657, 658, 658, 687, 687, 688, 688, 689, 689, 690, 690, 691, 691, 692, 692, 693, 693, 694, 694, 695, 695, 696, 696, 697, 697, 698, 698, 699, 699, 700, 700, 701, 701, 702, 702, 707, 707, 708, 708, 709, 709, 710, 710, 723, 723, 724, 724, 725, 725, 726, 726, 727, 727, 728, 728, 729, 729, 730, 730, 735, 735, 736, 736, 737, 737, 738, 738, 747, 747, 748, 748, 749, 749, 750, 750, 767, 767, 768, 768, 769, 769, 770, 770, 799, 799, 800, 800, 801, 801, 802, 802, 803, 803, 804, 804, 805, 805, 806, 806, 815, 815, 816, 816, 817, 817, 818, 818, 819, 819, 820, 820, 821, 821, 822, 822, 831, 831, 832, 832, 833, 833, 834, 834, 855, 855, 856, 856, 857, 857, 858, 858, 859, 859, 860, 860, 861, 861, 862, 862, 911, 911, 912, 912, 913, 913, 914, 914, 915, 915, 916, 916, 917, 917, 918, 918, 927, 927, 928, 928, 929, 929, 930, 930, 931, 931, 932, 932, 933, 933, 934, 934, 943, 943, 944, 944, 945, 945, 946, 946, 947, 947, 948, 948, 949, 949, 950, 950)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 2, 3, 4, 5, 6, 7, 8, 8, 7, 6, 7, 7, 8, 8, 9, 9, 5, 6, 7, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 8, 7, 4, 5, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 9, 9, 8, 9, 9, 7, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 9, 9, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 3, 4, 5, 6, 7, 8, 9, 9, 8, 7, 6, 5, 6, 6, 7, 8, 8, 9, 9, 7, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 5, 6, 7, 8, 8, 7, 6, 7, 8, 9, 9, 8, 7, 2, 3, 4, 5, 6, 7, 7, 8, 8, 9, 9, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 5, 6, 7, 7, 6, 4, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 6, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 8, 8, 9, 9, 6, 5, 6, 6, 7, 8, 8, 7, 8, 8, 9, 9, 4, 5, 6, 7, 7, 6, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 9, 9, 8, 1, 2, 3, 4, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 8, 9, 9, 5, 6, 7, 7, 8, 8, 9, 9, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 4, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 9, 9, 5, 6, 7, 8, 8, 9, 9, 7, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 3, 4, 5, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 6, 5, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 4, 5, 6, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 9, 9, 5, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 8, 7, 2, 3, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 8, 9, 9, 8, 5, 6, 7, 8, 8, 7, 8, 9, 9, 8, 6, 7, 8, 9, 9, 8, 7, 8, 8, 9, 9, 4, 5, 6, 7, 8, 8, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 8, 9, 9, 7, 8, 8, 5, 6, 7, 7, 6, 7, 7, 8, 8, 9, 9, 3, 4, 5, 6, 6, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 6, 7, 7, 8, 8, 4, 5, 6, 6, 7, 8, 9, 9, 8, 7, 5, 6, 6, 7, 7, 8, 9, 9, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 7, 7, 7, 7, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 9, 9, 7, 7, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 9, 8, 7, 8, 8, 6, 7, 8, 9, 9, 8, 7, 8, 8, 9, 9, 5, 6, 7, 8, 8, 9, 9, 7, 8, 8, 6, 7, 8, 8, 7, 4, 5, 6, 7, 8, 9, 9, 8, 7, 6, 7, 7, 8, 9, 9, 8, 5, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 6, 7, 8, 9, 9, 8, 7, 3, 4, 5, 6, 6, 7, 7, 8, 9, 9, 8, 9, 9, 5, 6, 7, 8, 9, 9, 8, 7, 6, 7, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 9, 9, 5, 6, 6, 7, 7, 8, 8, 9, 9, 2, 3, 4, 5, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 5, 6, 7, 7, 8, 8, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 9, 9, 4, 5, 6, 6, 7, 7, 8, 9, 9, 8, 5, 6, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 3, 4, 5, 6, 7, 8, 8, 7, 6, 7, 7, 8, 9, 9, 8, 9, 9, 5, 4, 5, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 6, 1, 2, 3, 4, 5, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 6, 7, 7, 8, 8, 9, 9, 5, 6, 7, 8, 9, 9, 8, 7, 8, 8, 9, 9, 6, 7, 8, 8, 7, 8, 8, 9, 9, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 9, 9, 8, 7, 8, 8, 9, 9, 5, 6, 7, 8, 8, 9, 9, 7, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 3, 4, 4, 5, 6, 7, 8, 8, 9, 9, 7, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 9, 9, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 2, 3, 4, 5, 5, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 9, 9, 4, 5, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 6, 7, 7, 8, 9, 9, 8, 9, 9, 5, 6, 7, 8, 8, 9, 9, 7, 6, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 4, 5, 6, 7, 8, 9, 9, 8, 7, 8, 8, 6, 5, 6, 7, 8, 8, 9, 9, 7, 8, 8, 6, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 6, 6, 6, 6, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 5, 5, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 6, 6, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 6, 6, 6, 6, 9, 9, 9, 9, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 2, 3, 4, 5, 6, 7, 7, 8, 9, 9, 8, 9, 9, 6, 7, 7, 5, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 6, 7, 7, 8, 8, 4, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 5, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 6, 7, 8, 9, 9, 8, 9, 9, 7, 3, 4, 5, 6, 6, 5, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 9, 9, 4, 5, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 2, 3, 4, 5, 6, 6, 7, 7, 8, 8, 9, 9, 5, 6, 7, 8, 9, 9, 8, 7, 8, 8, 6, 4, 5, 6, 7, 8, 9, 9, 8, 7, 6, 7, 7, 8, 8, 9, 9, 5, 6, 7, 8, 8, 9, 9, 7, 6, 3, 4, 5, 6, 6, 7, 7, 8, 9, 9, 8, 9, 9, 5, 6, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 9, 9, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 9, 9, 8, 7, 5, 6, 6, 7, 8, 8, 7, 1, 2, 3, 4, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 6, 7, 8, 8, 9, 9, 7, 5, 6, 7, 8, 8, 9, 9, 7, 6, 7, 8, 8, 9, 9, 7, 8, 8, 9, 9, 4, 5, 5, 6, 7, 7, 6, 7, 8, 9, 9, 8, 7, 8, 9, 9, 8, 3, 4, 5, 6, 7, 8, 9, 9, 8, 7, 6, 7, 8, 8, 7, 8, 9, 9, 8, 9, 9, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 9, 9, 8, 9, 9, 4, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 8, 9, 9, 6, 7, 8, 9, 9, 8, 7, 8, 8, 5, 6, 7, 7, 6, 2, 3, 4, 5, 5, 6, 7, 8, 8, 9, 9, 7, 6, 7, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 9, 9, 8, 9, 9, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 5, 6, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 3, 4, 5, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 8, 9, 9, 8, 9, 9, 6, 7, 7, 8, 8, 9, 9, 4, 5, 6, 7, 8, 8, 7, 6, 5, 6, 7, 8, 9, 9, 8, 9, 9, 7, 6, 7, 8, 9, 9, 8, 7, 8, 8, 9, 9, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 7, 7, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 7, 7, 7, 7, 8, 8, 7, 7, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 6, 6, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 6, 6, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 6, 6, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((16, 17, 23, 24, 26, 27, 39, 40, 43, 44, 46, 47, 51, 52, 54, 55, 61, 62, 64, 65, 69, 70, 74, 75, 77, 78, 81, 82, 84, 85, 92, 93, 103, 104, 116, 117, 121, 122, 133, 134, 146, 147, 152, 153, 157, 158, 169, 170, 172, 173, 180, 181, 183, 184, 197, 198, 209, 210, 227, 228, 245, 246, 253, 254, 259, 260, 263, 264, 271, 272, 274, 275, 278, 279, 284, 285, 289, 290, 292, 293, 299, 300, 306, 307, 310, 311, 313, 314, 322, 323, 327, 328, 334, 335, 339, 340, 342, 343, 347, 348, 350, 351, 354, 355, 363, 364, 366, 367, 371, 372, 378, 379, 382, 383, 385, 386, 407, 408, 417, 418, 423, 424, 429, 430, 439, 440, 442, 443, 448, 449, 462, 463, 473, 474, 476, 477, 492, 493, 502, 503, 505, 506, 507, 508, 513, 514, 517, 518, 519, 520, 523, 524, 527, 528, 529, 530, 537, 538, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 557, 558, 563, 564, 565, 566, 567, 568, 587, 588, 593, 594, 595, 596, 597, 598, 607, 608, 609, 610, 613, 614, 617, 618, 619, 620, 623, 624, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 641, 642, 643, 644, 645, 646, 649, 650, 651, 652, 655, 656, 657, 658, 659, 660, 661, 662, 665, 666, 667, 668, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 703, 704, 709, 710, 711, 712, 715, 716, 717, 718, 721, 722, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 763, 764, 765, 766, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 795, 796, 797, 798, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 827, 828, 829, 830, 831, 832, 833, 834, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 899, 900, 901, 902, 907, 908, 909, 910, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (9, 10, 18, 19, 24, 25, 31, 32, 46, 47, 54, 55, 61, 62, 66, 67, 72, 73, 84, 85, 87, 88, 93, 94, 112, 113, 117, 118, 120, 121, 129, 130, 139, 140, 144, 145, 149, 150, 152, 153, 166, 167, 169, 170, 174, 175, 183, 184, 192, 193, 196, 197, 211, 212, 214, 215, 223, 224, 226, 227, 230, 231, 243, 244, 248, 249, 255, 256, 261, 262, 267, 268, 276, 277, 288, 289, 294, 295, 301, 302, 308, 309, 313, 314, 323, 324, 329, 330, 332, 333, 337, 338, 343, 344, 346, 347, 350, 351, 357, 358, 361, 362, 364, 365, 375, 376, 379, 380, 385, 386, 390, 391, 393, 394, 400, 401, 405, 406, 412, 413, 415, 416, 422, 423, 443, 444, 446, 447, 450, 451, 453, 454, 459, 460, 463, 464, 466, 467, 473, 474, 485, 486, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 513, 514, 519, 520, 521, 522, 523, 524, 525, 526, 533, 534, 539, 540, 541, 542, 543, 544, 545, 546, 549, 550, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 567, 568, 569, 570, 571, 572, 577, 578, 581, 582, 583, 584, 585, 586, 587, 588, 597, 598, 601, 602, 603, 604, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 633, 634, 635, 636, 639, 640, 643, 644, 645, 646, 647, 648, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 663, 664, 669, 670, 671, 672, 673, 674, 675, 676, 681, 682, 683, 684, 685, 686, 687, 688, 691, 692, 693, 694, 695, 696, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 739, 740, 741, 742, 743, 744, 745, 746, 751, 752, 753, 754, 759, 760, 761, 762, 763, 764, 765, 766, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 795, 796, 797, 798, 803, 804, 805, 806, 807, 808, 809, 810, 815, 816, 817, 818, 819, 820, 821, 822, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 879, 880, 881, 882, 883, 884, 885, 886, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (10, 11, 13, 14, 23, 24, 28, 29, 40, 41, 43, 44, 50, 51, 55, 56, 61, 62, 66, 67, 72, 73, 75, 76, 87, 88, 92, 93, 95, 96, 100, 101, 105, 106, 108, 109, 116, 117, 119, 120, 123, 124, 126, 127, 131, 132, 134, 135, 138, 139, 141, 142, 153, 154, 159, 160, 171, 172, 180, 181, 187, 188, 199, 200, 202, 203, 209, 210, 212, 213, 217, 218, 229, 230, 248, 249, 251, 252, 258, 259, 266, 267, 273, 274, 278, 279, 289, 290, 294, 295, 303, 304, 313, 314, 316, 317, 328, 329, 331, 332, 338, 339, 341, 342, 346, 347, 351, 352, 371, 372, 387, 388, 390, 391, 395, 396, 398, 399, 402, 403, 405, 406, 412, 413, 415, 416, 419, 420, 422, 423, 431, 432, 434, 435, 438, 439, 441, 442, 448, 449, 462, 463, 465, 466, 471, 472, 477, 478, 485, 486, 487, 488, 491, 492, 493, 494, 497, 498, 499, 500, 501, 502, 503, 504, 511, 512, 513, 514, 521, 522, 523, 524, 525, 526, 527, 528, 531, 532, 537, 538, 539, 540, 551, 552, 555, 556, 557, 558, 559, 560, 565, 566, 567, 568, 573, 574, 577, 578, 581, 582, 583, 584, 591, 592, 593, 594, 595, 596, 599, 600, 601, 602, 605, 606, 607, 608, 611, 612, 613, 614, 615, 616, 617, 618, 627, 628, 633, 634, 635, 636, 637, 638, 639, 640, 647, 648, 649, 650, 651, 652, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 703, 704, 705, 706, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 731, 732, 733, 734, 739, 740, 741, 742, 743, 744, 745, 746, 751, 752, 753, 754, 755, 756, 757, 758, 759, 760, 761, 762, 763, 764, 765, 766, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 807, 808, 809, 810, 811, 812, 813, 814, 823, 824, 825, 826, 827, 828, 829, 830, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 863, 864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 919, 920, 921, 922, 923, 924, 925, 926, 935, 936, 937, 938, 939, 940, 941, 942, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
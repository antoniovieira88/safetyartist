
    -------------------------------------------------------------------
    -- File   : stimulus_list_distance
    -------------------------------------------------------------------
    -- Description : Synchronous 128 x 24 ROM.
    -------------------------------------------------------------------
    -- Revision:
    --     Date        Rev     Author                      Description
    --     12/07/2023  1.0     Henrique Lefundes da Silva  Creation.
    -------------------------------------------------------------------
    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    entity stimulus_list_distance is
    port (
            address   : in  std_logic_vector(6 downto 0);
            clk       : in  std_logic;
            out_rom   : out std_logic_vector(23 downto 0)
        );
    end entity stimulus_list_distance;
    
    -- Initial data explicitly declared
    architecture stimulus_list_distance_arch of stimulus_list_distance is
      type memory_struct is array(0 to 127) of std_logic_vector(23 downto 0);
    
    signal memory : memory_struct := ("000000100111110100000111",
 	 	 	 	"000000101000100110110001",
 	 	 	 	"000000101000010010101001",
 	 	 	 	"000000101010011111010101",
 	 	 	 	"000000101001011111100000",
 	 	 	 	"000000101000001010110000",
 	 	 	 	"000000100100110000101000",
 	 	 	 	"000000101011001100111011",
 	 	 	 	"000000101000100110110001",
 	 	 	 	"000000101000001010110000",
 	 	 	 	"000000100111110010101000",
 	 	 	 	"000000101001011011101001",
 	 	 	 	"000000100111110000110110",
 	 	 	 	"000000101000001100111001",
 	 	 	 	"000000101000010100110100",
 	 	 	 	"000000100111111101111001",
 	 	 	 	"000000100101101001000010",
 	 	 	 	"000000101000000010000010",
 	 	 	 	"000000100111101001001000",
 	 	 	 	"000000101010011110110011",
 	 	 	 	"000000100110011000100111",
 	 	 	 	"000000101001010100101001",
 	 	 	 	"000000100111000001101110",
 	 	 	 	"000000101000001010110000",
 	 	 	 	"000000101000110010010001",
 	 	 	 	"000000101011001100111011",
 	 	 	 	"000000101011000001010110",
 	 	 	 	"000000101001011111100000",
 	 	 	 	"000000101011001100111011",
 	 	 	 	"000000100100110000101000",
 	 	 	 	"000000101001011111100000",
 	 	 	 	"000000101000011110111101",
 	 	 	 	"000000101000010100101010",
 	 	 	 	"000000101011000001010110",
 	 	 	 	"000000101001001110001111",
 	 	 	 	"000000101001100100001101",
 	 	 	 	"000000100111011010000011",
 	 	 	 	"000000100111110111110011",
 	 	 	 	"000000101011001111010111",
 	 	 	 	"000000101000100010100100",
 	 	 	 	"000000101000001010110000",
 	 	 	 	"000000101000000010000010",
 	 	 	 	"000000100111001001111100",
 	 	 	 	"000000100111011110011110",
 	 	 	 	"000000100111110010101000",
 	 	 	 	"000000100111001000110100",
 	 	 	 	"000000101001010110000101",
 	 	 	 	"000000101000101001110111",
 	 	 	 	"000000100101010100010010",
 	 	 	 	"000000101011001111010111",
 	 	 	 	"000000101000110010010001",
 	 	 	 	"000000101001100101001000",
 	 	 	 	"000000101010011111010111",
 	 	 	 	"000000100111011110100110",
 	 	 	 	"000000100111011110100110",
 	 	 	 	"000000101001010100101001",
 	 	 	 	"000000101001100101001000",
 	 	 	 	"000000101000100010100100",
 	 	 	 	"000000100110101100100000",
 	 	 	 	"000000101000010010101001",
 	 	 	 	"000000100111110111110011",
 	 	 	 	"000000100111101001001000",
 	 	 	 	"000000100111001001111100",
 	 	 	 	"000000101011001111010111",
 	 	 	 	"000000100111110100000111",
 	 	 	 	"000000100110111001011001",
 	 	 	 	"000000101010011111010111",
 	 	 	 	"000000101000111101001110",
 	 	 	 	"000000101001101101111010",
 	 	 	 	"000000101000010010101001",
 	 	 	 	"000000101000010000100111",
 	 	 	 	"000000100111110000100011",
 	 	 	 	"000000100111110111110011",
 	 	 	 	"000000101001010110000101",
 	 	 	 	"000000101001011010010000",
 	 	 	 	"000000100101100110000100",
 	 	 	 	"000101011100001101101000",
 	 	 	 	"000101101010000001001011",
 	 	 	 	"000110101101101100111100",
 	 	 	 	"000110111011001111010111",
 	 	 	 	"000111101001000011101000",
 	 	 	 	"000111001100111010010111",
 	 	 	 	"000110100001100000110001",
 	 	 	 	"000101100110110100110111",
 	 	 	 	"000100010110111010110011",
 	 	 	 	"000010001001000001000110",
 	 	 	 	"000001111110110000101000",
 	 	 	 	"000101001101001011100010",
 	 	 	 	"000101110000111100110000",
 	 	 	 	"001000011100111111001011",
 	 	 	 	"000100101101111011110100",
 	 	 	 	"000100101101111011110100",
 	 	 	 	"000100101101111011110100",
 	 	 	 	"000100101101111011110100",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000",
 	 	 	 	"000000000000000000000000");
  
    begin
    -- Reads ROM position at every rising edge of 'clk'.
    process (clk)
    begin
    if (clk'event and clk = '1') then
        out_rom <= memory(to_integer(unsigned(address)));
      end if;
    end process;

  end architecture stimulus_list_distance_arch;  
  
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((2, 2, 1, 0, 0, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, 0, -2, -2, 0, 0, 1, -2, -2, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, 0, 2, 0, 1, -2, -2, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, 1, 0, 0, -2, -2, 0, -2, -2, 2, 1, -2, -2, 1, -2, -2, 1, 1, 0, 2, 0, -2, -2, 0, -2, -2, 0, 2, -2, -2, 0, -2, -2, 2, 1, 0, -2, -2, 0, -2, -2, 1, 0, -2, -2, 1, -2, -2, 0, 0, 1, 2, -2, -2, 1, -2, -2, 0, -2, 0, -2, -2, 2, 1, 0, -2, -2, 0, -2, -2, 0, 0, -2, -2, 0, -2, -2, -2, -2),
                (2, 2, 0, 0, 1, 1, -2, -2, 1, -2, -2, 1, 0, -2, -2, 0, -2, -2, 1, 0, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 2, 0, 1, 0, -2, -2, 1, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 0, 0, -2, -2, 0, -2, -2, 1, 0, -2, -2, 0, -2, -2, 1, 0, 2, 1, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 1, 0, -2, -2, 2, -2, -2, 0, 0, -2, -2, 1, -2, -2, 1, 1, -2, 0, 0, -2, -2, 1, -2, -2, 2, 1, 1, -2, -2, 0, -2, -2, 0, 0, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 2, 1, 1, 0, -2, -2, 1, -2, -2, 1, 1, -2, -2, -2, 2, 2, 0, -2, -2, 1, -2, -2, 0, 0, -2, -2, 0, -2, -2, 0, 1, 1, 0, -2, -2, 1, -2, -2, 0, 2, -2, -2, 1, -2, -2, 2, 1, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 2, 2, 1, 0, 1, -2, -2, 0, -2, -2, 1, 1, -2, -2, 0, -2, -2, 0, 1, 1, -2, -2, 0, -2, -2, 1, 1, -2, -2, 1, -2, -2, 2, 1, 1, 0, -2, -2, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, 2, 1, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, 1, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((134, 92, 2452, 20555, 11497, 850, -256, -256, 1445, -256, -256, 33658, 33480, -256, -256, 39875, -256, -256, 71611, 52468, 2580, -256, -256, 3044, -256, -256, 3440, 78159, -256, -256, 3441, -256, -256, 34515, 109, 16401, 1111, -256, -256, 2016, -256, -256, 1664, 5753, -256, -256, 2194, -256, -256, 3047, 47219, 47191, -256, -256, 53771, -256, -256, 109, 3048, -256, -256, 3650, -256, -256, 2261, 1141, 4962, 164, 1239, -256, -256, 2540, -256, -256, 6436, 164, -256, -256, 8005, -256, -256, 164, 1150, 15404, -256, -256, 13729, -256, -256, 1733, 11649, -256, -256, 1733, -256, -256, 39733, 27064, 2330, 164, -256, -256, 2434, -256, -256, 27500, -256, 29629, -256, -256, 164, 3354, 43199, -256, -256, 53938, -256, -256, 45425, 44970, -256, -256, 45941, -256, -256, -256, -256),
                (134, 92, 46435, 21468, 1120, 858, -256, -256, 1372, -256, -256, 1970, 24380, -256, -256, 38324, -256, -256, 3061, 60475, 2732, -256, -256, 67878, -256, -256, 81972, 3256, -256, -256, 88188, -256, -256, 109, 41144, 1755, 10120, -256, -256, 2240, -256, -256, 65357, 3023, -256, -256, 3330, -256, -256, 40626, 10008, 4736, -256, -256, 24412, -256, -256, 3039, 44924, -256, -256, 60228, -256, -256, 2204, 10292, 164, 881, 4387, -256, -256, 7834, -256, -256, 2683, 480, -256, -256, 834, -256, -256, 15589, 1529, 12856, -256, -256, 164, -256, -256, 21828, 21819, -256, -256, 2134, -256, -256, 3070, 2204, -256, 31703, 26991, -256, -256, 2716, -256, -256, 164, 3739, 3071, -256, -256, 67143, -256, -256, 44808, 36810, -256, -256, 3510, -256, -256, -256, -256, -256, -256, -256, -256),
                (37372, 1678, 92, 1370, 593, 2543, -256, -256, 599, -256, -256, 1675, 1531, -256, -256, -256, 134, 109, 10418, -256, -256, 712, -256, -256, 6429, 2683, -256, -256, 11430, -256, -256, 24695, 1857, 1819, 16620, -256, -256, 1843, -256, -256, 21790, 164, -256, -256, 2200, -256, -256, 134, 2170, 28137, -256, -256, 35847, -256, -256, 30576, 2453, -256, -256, 30758, -256, -256, 109, 92, 2741, 49884, 2332, -256, -256, 52303, -256, -256, 3125, 2742, -256, -256, 83281, -256, -256, 56195, 2692, 2414, -256, -256, 52811, -256, -256, 3269, 3132, -256, -256, 3270, -256, -256, 134, 3011, 2824, 38227, -256, -256, 2824, -256, -256, 3013, 87008, -256, -256, 3567, -256, -256, 164, 3383, 3034, -256, -256, 3393, -256, -256, 42299, 42279, -256, -256, 3438, -256, -256, -256, -256)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((38, 38, 37, 40, 18, 11, 34, 0, 26, 41, 0, 42, 33, 33, 0, 43, 40, 43, 32, 5, 0, 3, 0, 17, 34, 0, 42, 42, 35, 43, 39, 0, 39, 38, 16, 16, 10, 30, 1, 22, 40, 2, 17, 32, 9, 38, 3, 12, 0, 42, 42, 38, 38, 0, 43, 41, 43, 37, 36, 0, 36, 38, 38, 33, 39, 41, 42, 12, 14, 0, 23, 9, 3, 22, 43, 29, 28, 29, 43, 42, 43, 40, 40, 33, 0, 43, 40, 2, 42, 40, 41, 1, 43, 40, 0, 40, 36, 4, 0, 2, 2, 2, 0, 1, 0, 14, 43, 14, 6, 16, 42, 42, 42, 28, 43, 39, 1, 43, 42, 34, 35, 0, 43, 39, 43, 43, 43),
                (38, 38, 37, 18, 10, 31, 34, 22, 1, 13, 0, 25, 41, 34, 42, 4, 1, 10, 41, 42, 39, 42, 9, 43, 42, 43, 35, 4, 9, 1, 42, 33, 43, 38, 38, 18, 34, 13, 41, 4, 13, 0, 42, 35, 41, 2, 43, 43, 41, 38, 19, 7, 3, 10, 23, 18, 27, 42, 43, 40, 43, 39, 7, 42, 39, 41, 13, 11, 28, 13, 43, 1, 0, 5, 15, 2, 11, 0, 21, 41, 6, 42, 32, 42, 40, 43, 3, 2, 5, 43, 39, 39, 0, 43, 43, 43, 36, 37, 0, 37, 3, 1, 16, 42, 43, 42, 35, 34, 34, 0, 34, 20, 0, 43, 35, 2, 0, 11, 43, 43, 42, 0, 0, 0, 0, 0, 0),
                (38, 19, 34, 32, 35, 40, 8, 43, 31, 0, 31, 17, 16, 20, 10, 43, 35, 34, 34, 16, 41, 34, 39, 30, 36, 12, 4, 21, 41, 32, 42, 5, 1, 8, 9, 1, 27, 5, 2, 15, 1, 0, 0, 1, 4, 18, 0, 14, 9, 36, 23, 40, 1, 1, 5, 21, 17, 40, 2, 25, 32, 24, 42, 41, 41, 42, 38, 43, 4, 43, 41, 43, 36, 38, 0, 38, 34, 2, 42, 41, 32, 42, 43, 33, 4, 2, 15, 42, 43, 43, 42, 40, 0, 40, 42, 42, 43, 43, 37, 43, 41, 0, 41, 38, 9, 0, 43, 38, 39, 35, 42, 42, 42, 43, 41, 39, 32, 39, 42, 37, 37, 0, 43, 43, 42, 43, 43)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 3, 4, 5, 6, -1, -1, 9, -1, -1, 12, 13, -1, -1, 16, -1, -1, 19, 20, 21, -1, -1, 24, -1, -1, 27, 28, -1, -1, 31, -1, -1, 34, 35, 36, 37, -1, -1, 40, -1, -1, 43, 44, -1, -1, 47, -1, -1, 50, 51, 52, -1, -1, 55, -1, -1, 58, 59, -1, -1, 62, -1, -1, 65, 66, 67, 68, 69, -1, -1, 72, -1, -1, 75, 76, -1, -1, 79, -1, -1, 82, 83, 84, -1, -1, 87, -1, -1, 90, 91, -1, -1, 94, -1, -1, 97, 98, 99, 100, -1, -1, 103, -1, -1, 106, 125, 108, -1, -1, 111, 112, 113, -1, -1, 116, -1, -1, 119, 120, -1, -1, 123, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, -1, -1, 9, -1, -1, 12, 13, -1, -1, 16, -1, -1, 19, 20, 21, -1, -1, 24, -1, -1, 27, 28, -1, -1, 31, -1, -1, 34, 35, 36, 37, -1, -1, 40, -1, -1, 43, 44, -1, -1, 47, -1, -1, 50, 51, 52, -1, -1, 55, -1, -1, 58, 59, -1, -1, 62, -1, -1, 65, 66, 67, 68, 69, -1, -1, 72, -1, -1, 75, 76, -1, -1, 79, -1, -1, 82, 83, 84, -1, -1, 87, -1, -1, 90, 91, -1, -1, 94, -1, -1, 97, 98, 121, 100, 101, -1, -1, 104, -1, -1, 107, 108, 109, -1, -1, 112, -1, -1, 115, 116, -1, -1, 119, -1, -1, 123, 125, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, -1, -1, 9, -1, -1, 12, 13, -1, -1, 125, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1, 32, 33, 34, 35, -1, -1, 38, -1, -1, 41, 42, -1, -1, 45, -1, -1, 48, 49, 50, -1, -1, 53, -1, -1, 56, 57, -1, -1, 60, -1, -1, 63, 64, 65, 66, 67, -1, -1, 70, -1, -1, 73, 74, -1, -1, 77, -1, -1, 80, 81, 82, -1, -1, 85, -1, -1, 88, 89, -1, -1, 92, -1, -1, 95, 96, 97, 98, -1, -1, 101, -1, -1, 104, 105, -1, -1, 108, -1, -1, 111, 112, 113, -1, -1, 116, -1, -1, 119, 120, -1, -1, 123, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((64, 33, 18, 11, 8, 7, -1, -1, 10, -1, -1, 15, 14, -1, -1, 17, -1, -1, 26, 23, 22, -1, -1, 25, -1, -1, 30, 29, -1, -1, 32, -1, -1, 49, 42, 39, 38, -1, -1, 41, -1, -1, 46, 45, -1, -1, 48, -1, -1, 57, 54, 53, -1, -1, 56, -1, -1, 61, 60, -1, -1, 63, -1, -1, 96, 81, 74, 71, 70, -1, -1, 73, -1, -1, 78, 77, -1, -1, 80, -1, -1, 89, 86, 85, -1, -1, 88, -1, -1, 93, 92, -1, -1, 95, -1, -1, 110, 105, 102, 101, -1, -1, 104, -1, -1, 107, 126, 109, -1, -1, 118, 115, 114, -1, -1, 117, -1, -1, 122, 121, -1, -1, 124, -1, -1, -1, -1),
                (64, 33, 18, 11, 8, 7, -1, -1, 10, -1, -1, 15, 14, -1, -1, 17, -1, -1, 26, 23, 22, -1, -1, 25, -1, -1, 30, 29, -1, -1, 32, -1, -1, 49, 42, 39, 38, -1, -1, 41, -1, -1, 46, 45, -1, -1, 48, -1, -1, 57, 54, 53, -1, -1, 56, -1, -1, 61, 60, -1, -1, 63, -1, -1, 96, 81, 74, 71, 70, -1, -1, 73, -1, -1, 78, 77, -1, -1, 80, -1, -1, 89, 86, 85, -1, -1, 88, -1, -1, 93, 92, -1, -1, 95, -1, -1, 106, 99, 122, 103, 102, -1, -1, 105, -1, -1, 114, 111, 110, -1, -1, 113, -1, -1, 118, 117, -1, -1, 120, -1, -1, 124, 126, -1, -1, -1, -1),
                (62, 31, 16, 11, 8, 7, -1, -1, 10, -1, -1, 15, 14, -1, -1, 126, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1, 47, 40, 37, 36, -1, -1, 39, -1, -1, 44, 43, -1, -1, 46, -1, -1, 55, 52, 51, -1, -1, 54, -1, -1, 59, 58, -1, -1, 61, -1, -1, 94, 79, 72, 69, 68, -1, -1, 71, -1, -1, 76, 75, -1, -1, 78, -1, -1, 87, 84, 83, -1, -1, 86, -1, -1, 91, 90, -1, -1, 93, -1, -1, 110, 103, 100, 99, -1, -1, 102, -1, -1, 107, 106, -1, -1, 109, -1, -1, 118, 115, 114, -1, -1, 117, -1, -1, 122, 121, -1, -1, 124, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 1, 2, 3, 4, 5, 5, 4, 8, 8, 3, 11, 12, 12, 11, 15, 15, 2, 18, 19, 20, 20, 19, 23, 23, 18, 26, 27, 27, 26, 30, 30, 1, 33, 34, 35, 36, 36, 35, 39, 39, 34, 42, 43, 43, 42, 46, 46, 33, 49, 50, 51, 51, 50, 54, 54, 49, 57, 58, 58, 57, 61, 61, 0, 64, 65, 66, 67, 68, 68, 67, 71, 71, 66, 74, 75, 75, 74, 78, 78, 65, 81, 82, 83, 83, 82, 86, 86, 81, 89, 90, 90, 89, 93, 93, 64, 96, 97, 98, 99, 99, 98, 102, 102, 97, 105, 105, 107, 107, 96, 110, 111, 112, 112, 111, 115, 115, 110, 118, 119, 119, 118, 122, 122, 106, 106),
                (-1, 0, 1, 2, 3, 4, 5, 5, 4, 8, 8, 3, 11, 12, 12, 11, 15, 15, 2, 18, 19, 20, 20, 19, 23, 23, 18, 26, 27, 27, 26, 30, 30, 1, 33, 34, 35, 36, 36, 35, 39, 39, 34, 42, 43, 43, 42, 46, 46, 33, 49, 50, 51, 51, 50, 54, 54, 49, 57, 58, 58, 57, 61, 61, 0, 64, 65, 66, 67, 68, 68, 67, 71, 71, 66, 74, 75, 75, 74, 78, 78, 65, 81, 82, 83, 83, 82, 86, 86, 81, 89, 90, 90, 89, 93, 93, 64, 96, 97, 97, 99, 100, 100, 99, 103, 103, 96, 106, 107, 108, 108, 107, 111, 111, 106, 114, 115, 115, 114, 118, 118, 98, 98, 121, 121, 122, 122),
                (-1, 0, 1, 2, 3, 4, 5, 5, 4, 8, 8, 3, 11, 12, 12, 11, 2, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28, 1, 31, 32, 33, 34, 34, 33, 37, 37, 32, 40, 41, 41, 40, 44, 44, 31, 47, 48, 49, 49, 48, 52, 52, 47, 55, 56, 56, 55, 59, 59, 0, 62, 63, 64, 65, 66, 66, 65, 69, 69, 64, 72, 73, 73, 72, 76, 76, 63, 79, 80, 81, 81, 80, 84, 84, 79, 87, 88, 88, 87, 91, 91, 62, 94, 95, 96, 97, 97, 96, 100, 100, 95, 103, 104, 104, 103, 107, 107, 94, 110, 111, 112, 112, 111, 115, 115, 110, 118, 119, 119, 118, 122, 122, 15, 15)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 1, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 6, 6),
                (0, 1, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 1, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 2, 3, 4, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 5, 5, 6, 6, 6, 6),
                (0, 1, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 1, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 2, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 3, 4, 5, 6, 6, 5, 6, 6, 4, 5, 6, 6, 5, 6, 6, 6, 6)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((6, 7, 9, 10, 13, 14, 16, 17, 21, 22, 24, 25, 28, 29, 31, 32, 37, 38, 40, 41, 44, 45, 47, 48, 52, 53, 55, 56, 59, 60, 62, 63, 69, 70, 72, 73, 76, 77, 79, 80, 84, 85, 87, 88, 91, 92, 94, 95, 100, 101, 103, 104, 108, 109, 113, 114, 116, 117, 120, 121, 123, 124, 125, 126),
                (6, 7, 9, 10, 13, 14, 16, 17, 21, 22, 24, 25, 28, 29, 31, 32, 37, 38, 40, 41, 44, 45, 47, 48, 52, 53, 55, 56, 59, 60, 62, 63, 69, 70, 72, 73, 76, 77, 79, 80, 84, 85, 87, 88, 91, 92, 94, 95, 101, 102, 104, 105, 109, 110, 112, 113, 116, 117, 119, 120, 123, 124, 125, 126),
                (6, 7, 9, 10, 13, 14, 19, 20, 22, 23, 26, 27, 29, 30, 35, 36, 38, 39, 42, 43, 45, 46, 50, 51, 53, 54, 57, 58, 60, 61, 67, 68, 70, 71, 74, 75, 77, 78, 82, 83, 85, 86, 89, 90, 92, 93, 98, 99, 101, 102, 105, 106, 108, 109, 113, 114, 116, 117, 120, 121, 123, 124, 125, 126)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 2, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 2, 1, 0, 1, 2, 2, 1, -2, 1, 1, 1, 1, 1, 1, 0, 0, 2, 2, 2, 0, -2, 0, 0, 0, 0, 2, -2, -2, 2, 0, -2, -2, 2, -2, 1, 0, 0, 0, 2, 0, 1, -2, -2, -2, 1, 1, 0, 2, -2, -2, 0, 1, -2, 0, 0, 0, -2, -2, -2, 0, -2, 1, 1, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, 2, -2, -2, 0, 0, -2, -2, -2, 1, 2, 0, 0, 0, 0, -2, -2, -2, -2, -2, -2, 2, 2, 2, -2, -2, -2, -2, -2, -2, 2, -2, -2, 1, -2, -2, -2, 2, -2, -2, -2, -2, 1, 1, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, 2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 2, 2, 0, 0, 2, 2, 1, 2, 0, 0, 0, 1, 1, 2, 1, -2, -2, -2, 1, 0, 1, 2, 0, 1, 1, 0, 1, 2, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, -2, -2, 1, 0, 0, 2, 1, 1, 2, 1, 0, 2, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2, 1, 1, -2, -2, 2, 0, 2, 0, 1, 0, -2, 1, -2, -2, 2, 0, 0, 1, 2, 1, 2, -2, 0, -2, -2, -2, 1, -2, -2, -2, 1, 1, 1, 0, 2, 1, -2, -2, 0, -2, 1, -2, -2, -2, 2, 1, 1, 1, 0, 1, -2, -2, 1, -2, 0, -2, -2, -2, -2, 2, -2, -2, 2, 2, -2, -2, 1, 1, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, 0, -2, -2, 0, 0, -2, -2, -2, -2, 1, 1, 1, 2, -2, 2, -2, -2, 1, -2, 0, 0, -2, -2, -2, -2, -2, 2, 0, -2, 0, -2, -2, 0, 2, -2, -2, -2, 1, -2, -2, -2, 0, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, 0, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 1, 1, 2, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, 1, -2, -2, -2, 0, 0, -2, -2, -2, 1, -2, -2, -2, 1, 1, -2, 2, 0, -2, -2, -2, 1, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 1, 2, 1, 2, 1, 1, -2, -2, 0, 0, 0, 1, -2, -2, 0, 0, 0, 0, -2, -2, 0, -2, -2, -2, 1, 0, -2, -2, -2, -2, 1, 1, 1, 2, 1, 0, 1, 1, -2, -2, 1, 1, -2, 2, -2, 2, 0, -2, -2, -2, -2, -2, -2, -2, 2, 0, -2, -2, -2, -2, -2, -2, 1, 1, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, 0, 0, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((1844779, 60500, 2787704, 525669, 931537, 33517, 49724, 731177, 86054, 93167, 118138, 90146, 3502, 1261392, 4285, 169601, 332826, 13873, 27573, 2299169, 2134159, 584219, 789669, 1511576, 1265664, 4285, 859141, 91164, 102030, 4285, 3502, 72202, 79676, 37598, 45252, 69268, 75834, 59449, 119402, 4285, 83297, 20389, 12197, 4285, 5238, 73530, -8192, 67338, 71920, 102609, 105000, 87816, 99065, 1398013, 1597045, 2929, 3502, 3502, 1764404, -8192, 1658101, 209818, 307657, 2494762, 2929, -8192, -8192, 2929, 2077459, -8192, -8192, 4285, -8192, 113471, 2481044, 705788, 582832, 4285, 328740, 105953, -8192, -8192, -8192, 103216, 110933, 1165428, 5238, -8192, -8192, 409771, 43279, -8192, 1066660, 2208278, 2011359, -8192, -8192, -8192, 2050314, -8192, 25471, 44629, -8192, -8192, -8192, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, 237255, -8192, -8192, -8192, -8192, -8192, 3502, -8192, -8192, 2909358, 644761, -8192, -8192, -8192, 54509, 2929, 446858, 449265, 735798, 825405, -8192, -8192, -8192, -8192, -8192, -8192, 5238, 4285, 2929, -8192, -8192, -8192, -8192, -8192, -8192, 4285, -8192, -8192, 55406, -8192, -8192, -8192, 3502, -8192, -8192, -8192, -8192, 62669, 23213, -8192, -8192, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, -8192, 87323, -8192, -8192, -8192, 55494, -8192, 5238, -8192, -8192, 812820, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 522747, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192),
                (1600214, 42280, 2333905, 329127, 1092678, 12601, 399681, 94614, 2785418, 85962, 4285, 60783, 76578, 70388, 88354, 2093067, 1750943, 61440, 244055, 39194, 79710, 615745, 829863, 490891, 771969, 83641, 2929, 1966510, 1712790, 4285, 5238, 1299388, 1098606, 4285, 2929, 66531, 2929, 1516226, 1114046, 194600, 30506, 28609, 4285, 53868, -8192, -8192, -8192, 35120, 430080, 31915, 4285, 1918343, 94274, 104611, 2831086, 102371, 2929, 106935, 3502, 98280, 3502, 99938, 118598, 93976, 100753, 1186963, 1478092, -8192, -8192, 108586, 1778010, 450727, 5238, 47860, 60293, 2929, 107039, 1607436, 5238, 77362, 3502, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 53926, 60255, -8192, -8192, 3502, 345973, 3502, 1756569, 87575, 1606175, -8192, 34974, -8192, -8192, 3502, 1145598, 736353, 73174, 4285, 83146, 3502, -8192, 1265724, -8192, -8192, -8192, 115080, -8192, -8192, -8192, 18368, 27533, 23023, 194667, 5238, 84872, -8192, -8192, 2480643, -8192, 112870, -8192, -8192, -8192, 3502, 102894, 98245, 96722, 36116, 6987, -8192, -8192, 114336, -8192, 2142181, -8192, -8192, -8192, -8192, 2929, -8192, -8192, 4285, 4285, -8192, -8192, 105501, 105884, 98108, 2929, 2474345, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 121528, 140595, -8192, -8192, 1796580, 1926189, -8192, -8192, -8192, -8192, 39219, 42205, 37404, 4285, -8192, 2929, -8192, -8192, 40221, -8192, 403566, 451085, -8192, -8192, -8192, -8192, -8192, 2929, 1788969, -8192, 1643283, -8192, -8192, 1149787, 2929, -8192, -8192, -8192, 10256, -8192, -8192, -8192, 2680321, 110737, 106863, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 3502, 2012636, -8192, -8192, -8192, 86839, -8192, -8192, -8192, 39139, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 1751766, -8192, -8192, -8192, 61298, 74331, 5238, -8192, -8192, -8192, -8192, -8192, -8192, 3236, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 40425, 42215, -8192, -8192, -8192, 2423576, 2418123, -8192, -8192, -8192, 110564, -8192, -8192, -8192, 110466, 117066, -8192, 2929, 2794312, -8192, -8192, -8192, 114933, -8192, -8192, -8192, -8192, 36529, -8192, -8192, -8192, -8192, -8192, -8192, 61291, 659498, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 520375, -8192, -8192, -8192, -8192, -8192, 117082, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192),
                (1881051, 39120, 2417815, 325473, 1142411, 15876, 397028, 67490, 78286, 69527, 4285, 95658, 2786086, 89411, 3502, 103605, 4285, 83279, 95145, -8192, -8192, 775038, 901648, 543896, 58925, -8192, -8192, 84591, 237589, 46910, 102020, -8192, -8192, 2054985, -8192, -8192, -8192, 68222, 1304821, -8192, -8192, -8192, -8192, 103920, 120411, 100064, 2929, 109474, 2450850, 19167, 28247, -8192, -8192, 32040, 38493, -8192, 4285, -8192, 2929, 2087171, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 2929, 2254823, -8192, -8192, -8192, -8192, -8192, -8192, 72785, 84541, -8192, -8192, -8192, -8192, -8192, 2514692, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 473308, -8192, -8192, 2878438, 3443625, -8192, -8192, -8192, -8192, 111008, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((1094, 521, 1348, 965, 200, 416, 1319, 19, 454, 1251, 1365, 1364, 863, 958, 195, 795, 96, 264, 1263, 483, 1283, 1363, 1136, 58, 465, 527, 1355, 92, 803, 631, 1207, 366, 1216, 9, 311, 2, 85, 704, 53, 319, 6, 145, 1329, 812, 57, 1015, 1365, 68, 1014, 225, 833, 3, 163, 1186, 474, 824, 101, 442, 12, 1365, 733, 1356, 965, 1272, 511, 198, 1064, 570, 39, 163, 1108, 1126, 1365, 180, 1138, 291, 1195, 542, 1346, 777, 1365, 522, 1365, 1328, 195, 482, 27, 379, 1157, 543, 1302, 1365, 919, 257, 1039, 910, 1342, 1365, 1303, 0, 195, 1316, 1365, 473, 1365, 140, 945, 1365, 975, 18, 294, 0, 1365, 69, 0, 433, 0, 614, 1365, 1189, 1365, 1365, 1336, 14, 0, 195, 1109, 159, 703, 14, 280, 1293, 634, 0, 396, 118, 993, 287, 1365, 3, 124, 1006, 1365, 759, 1365, 310, 1078, 0, 282, 0, 910, 780, 1365, 228, 1365, 162, 0, 455, 1365, 0, 488, 1278, 1365, 53, 735, 320, 24, 1143, 1365, 862, 1365, 210, 1024, 52, 0, 1365, 853, 759, 1365, 32, 0, 0, 216, 1365, 341, 53, 398, 256, 0, 0, 80, 0, 178, 1365, 1092, 0, 54, 0, 50, 1365, 248, 1365, 273, 0, 248, 1365, 1092, 0, 512, 420, 62, 1365, 1092, 0, 35, 1241, 1365, 0, 15, 0, 114, 910, 1326, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 228, 228, 1365, 1365, 0, 0, 455, 455, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 228, 228, 228, 228, 1365, 1365, 1365, 1365, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 455, 455, 455, 455, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365),
                (888, 255, 1302, 845, 117, 219, 1332, 955, 1357, 1308, 301, 52, 360, 1226, 129, 121, 1189, 713, 111, 100, 1345, 216, 16, 48, 979, 1362, 918, 322, 1250, 401, 61, 177, 1323, 654, 1231, 1349, 853, 231, 1217, 47, 480, 1291, 137, 411, 1365, 941, 105, 947, 1358, 1299, 260, 100, 1081, 1263, 1365, 1357, 691, 76, 1263, 51, 340, 177, 1232, 26, 307, 819, 112, 119, 1203, 768, 1357, 12, 281, 155, 1311, 768, 78, 1165, 319, 7, 335, 183, 1152, 303, 1365, 710, 77, 52, 910, 940, 1347, 1365, 439, 78, 1170, 875, 1347, 195, 1256, 0, 522, 1365, 218, 637, 1318, 4, 67, 377, 26, 137, 1365, 149, 1365, 0, 1195, 158, 1365, 59, 501, 21, 200, 1038, 33, 137, 3, 43, 1092, 1006, 1365, 455, 1365, 1138, 0, 223, 28, 65, 1170, 13, 372, 1365, 0, 1295, 0, 1179, 0, 1365, 735, 1365, 869, 0, 1365, 106, 10, 54, 423, 546, 1271, 1363, 1138, 171, 1365, 34, 455, 1365, 22, 1365, 0, 49, 1365, 0, 1308, 204, 11, 131, 5, 13, 1241, 55, 512, 1365, 228, 1365, 105, 1227, 1363, 1343, 341, 1365, 993, 0, 1365, 195, 1365, 5, 119, 1365, 91, 910, 1365, 1365, 1231, 735, 1365, 195, 1365, 1365, 1219, 546, 1365, 0, 1365, 975, 1365, 1365, 0, 287, 39, 161, 1365, 85, 1365, 910, 0, 1365, 1024, 1365, 975, 92, 10, 19, 585, 683, 1336, 1024, 1348, 0, 341, 683, 0, 0, 683, 683, 0, 683, 1365, 683, 0, 1365, 1062, 1365, 975, 1155, 1365, 1365, 0, 1, 28, 137, 0, 52, 1252, 0, 44, 1365, 1024, 0, 1365, 256, 0, 0, 152, 1365, 1195, 0, 71, 1364, 1170, 0, 1365, 1365, 1303, 1073, 1365, 1252, 0, 98, 0, 67, 1365, 1331, 1365, 1365, 745, 228, 1365, 1365, 0, 1195, 1365, 1365, 0, 0, 171, 1365, 0, 1, 40, 114, 0, 44, 1, 22, 1365, 0, 29, 37, 1, 1365, 1333, 975, 1365, 0, 9, 1365, 1356, 0, 1365, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 683, 683, 0, 0, 0, 0, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365),
                (750, 217, 1313, 803, 119, 188, 1341, 45, 365, 1251, 140, 952, 1356, 1339, 345, 80, 1047, 57, 413, 1132, 214, 148, 7, 53, 920, 1289, 545, 519, 78, 109, 1335, 15, 269, 671, 1365, 198, 1214, 1357, 968, 484, 1256, 388, 33, 1237, 1365, 1359, 593, 67, 1319, 30, 391, 1365, 112, 943, 1364, 1365, 228, 1365, 1021, 359, 1365, 94, 1214, 42, 503, 85, 1365, 221, 28, 53, 643, 175, 12, 910, 1365, 2, 33, 127, 4, 956, 1365, 1365, 1217, 910, 1365, 1365, 1209, 180, 16, 7, 88, 1365, 1280, 0, 1365, 1365, 1280, 683, 1365, 11, 1, 1354, 1365, 1365, 1124, 1132, 1132, 214, 214, 1289, 1289, 545, 545, 15, 15, 269, 269, 1365, 1365, 198, 198, 1214, 1214, 484, 484, 1256, 1256, 388, 388, 33, 33, 1365, 1365, 112, 112, 1365, 1365, 1365, 1365, 1365, 1365, 94, 94, 1214, 1214, 42, 42, 503, 503, 85, 85, 1365, 1365, 53, 53, 643, 643, 175, 175, 12, 12, 910, 910, 1365, 1365, 127, 127, 4, 4, 956, 956, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 1365, 1365, 1209, 1209, 180, 180, 16, 16, 7, 7, 88, 88, 1365, 1365, 0, 0, 1365, 1365, 683, 683, 1365, 1365, 11, 11, 1, 1, 1365, 1365, 1365, 1365, 1124, 1124, 1132, 1132, 1132, 1132, 214, 214, 214, 214, 1289, 1289, 1289, 1289, 545, 545, 545, 545, 15, 15, 15, 15, 269, 269, 269, 269, 1365, 1365, 1365, 1365, 198, 198, 198, 198, 1214, 1214, 1214, 1214, 484, 484, 484, 484, 1256, 1256, 1256, 1256, 388, 388, 388, 388, 33, 33, 33, 33, 1365, 1365, 1365, 1365, 112, 112, 112, 112, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 94, 94, 94, 94, 1214, 1214, 1214, 1214, 42, 42, 42, 42, 503, 503, 503, 503, 85, 85, 85, 85, 1365, 1365, 1365, 1365, 53, 53, 53, 53, 643, 643, 643, 643, 175, 175, 175, 175, 12, 12, 12, 12, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 127, 127, 127, 127, 4, 4, 4, 4, 956, 956, 956, 956, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1209, 1209, 1209, 1209, 180, 180, 180, 180, 16, 16, 16, 16, 7, 7, 7, 7, 88, 88, 88, 88, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 11, 11, 11, 11, 1, 1, 1, 1, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1124, 1124, 1124, 1124, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 683, 683, 683, 683, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 9, 5, 7, 15, 21, 35, 13, 11, 121, 97, 19, 29, 23, 17, 33, 37, 61, 49, 71, 101, 25, 51, 27, 75, 119, 85, 53, 31, 45, 55, 91, 113, 43, 123, 39, 41, 99, 47, 179, 133, 193, 89, 129, 59, 223, 155, 131, 67, 63, 173, 57, 95, 65, 87, 109, 69, 197, 225, 81, 161, 77, 167, 73, -1, -1, 93, 189, -1, -1, 79, 227, 187, 143, 127, 151, 145, 215, 83, 229, -1, -1, 211, 209, 125, 195, -1, -1, 105, 205, 231, 103, 135, 117, -1, -1, 233, 141, 235, 115, 107, 237, -1, -1, -1, -1, 239, 111, -1, -1, 241, 243, 147, 245, -1, -1, -1, -1, 177, 247, 249, 157, 139, 251, -1, -1, 165, 171, 213, 163, 221, 137, -1, -1, -1, -1, -1, -1, 217, 159, 153, 253, -1, -1, -1, -1, 255, 149, -1, -1, 183, 257, 259, 261, 185, 263, 265, 267, 269, 199, 175, 271, -1, -1, -1, -1, 169, 273, -1, -1, -1, -1, 203, 275, -1, -1, 201, 277, 181, 279, 281, 207, -1, -1, -1, -1, -1, -1, 283, 191, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 285, 219, -1, -1, -1, -1, 287, 289, -1, -1, 291, 293, 295, 297, -1, -1, 299, 301, -1, -1, 303, 305, 307, 309, -1, -1, -1, -1, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, -1, -1, -1, -1, 331, 333, 335, 337, -1, -1, 339, 341, 343, 345, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 347, 349, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 351, 353, 355, 357, -1, -1, -1, -1, 359, 361, 363, 365, 367, 369, 371, 373, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, -1, -1, -1, -1, -1, -1, -1, -1, 399, 401, 403, 405, 407, 409, 411, 413, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 415, 417, 419, 421, 423, 425, 427, 429, -1, -1, -1, -1, -1, -1, -1, -1, 431, 433, 435, 437, 439, 441, 443, 445, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 447, 449, 451, 453, 455, 457, 459, 461, 463, 465, 467, 469, 471, 473, 475, 477, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 11, 17, 47, 9, 53, 25, 15, 21, 13, 35, 29, 59, 69, 19, 39, 137, 211, 23, 105, 71, 33, 199, 27, 51, 95, 31, 63, 79, 231, 43, 89, 205, 37, 111, 103, 119, 41, 187, 99, 45, 327, -1, -1, 49, 183, 147, 93, 177, 143, 55, 289, 157, 57, 215, 127, 133, 61, 75, 141, 151, 65, 67, 87, -1, -1, 77, 297, 193, 73, 85, 165, 83, 171, 155, 115, 307, 81, -1, -1, -1, -1, -1, -1, -1, -1, 91, 223, -1, -1, 235, 243, 97, 251, 181, 169, 329, 101, -1, -1, 113, 233, 255, 107, 109, 123, 117, 331, 161, 333, -1, -1, 267, 335, -1, -1, 173, 121, 145, 163, 125, 315, -1, -1, 129, 337, 131, 339, -1, -1, 135, 227, 167, 249, 301, 139, 341, 343, 225, 345, 197, 347, -1, -1, 349, 149, 351, 353, 153, 261, -1, -1, 221, 247, 279, 159, 239, 355, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 175, 313, -1, -1, 269, 179, -1, -1, -1, -1, 185, 275, 263, 191, 357, 189, -1, -1, 241, 359, 305, 195, -1, -1, -1, -1, 361, 201, 203, 363, 245, 365, 367, 207, 209, 369, -1, -1, 213, 371, 373, 375, 217, 285, 219, 377, -1, -1, -1, -1, -1, -1, -1, -1, 229, 273, -1, -1, 379, 271, -1, -1, 381, 237, -1, -1, 383, 385, -1, -1, 387, 389, -1, -1, -1, -1, -1, -1, 253, 391, -1, -1, 309, 257, 259, 393, -1, -1, -1, -1, 395, 265, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 317, 277, 397, 399, 401, 281, 283, 403, -1, -1, 287, 405, -1, -1, 291, 323, 407, 293, 295, 409, 411, 413, 299, 415, 417, 419, 421, 303, -1, -1, -1, -1, -1, -1, 311, 321, -1, -1, -1, -1, -1, -1, 423, 319, -1, -1, -1, -1, 425, 325, 427, 429, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 431, 433, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 435, 437, -1, -1, -1, -1, 439, 441, -1, -1, -1, -1, 443, 445, 447, 449, -1, -1, 451, 453, -1, -1, 455, 457, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 459, 461, -1, -1, -1, -1, 463, 465, 467, 469, -1, -1, -1, -1, 471, 473, -1, -1, -1, -1, -1, -1, -1, -1, 475, 477, 479, 481, 483, 485, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 487, 489, 491, 493, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 495, 497, 499, 501, -1, -1, -1, -1, -1, -1, -1, -1, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 11, 5, 7, 27, 53, 21, 9, 37, 17, 13, 43, 57, 15, 67, 33, 41, 19, 105, 107, 23, 75, 31, 25, 109, 111, 29, 49, 63, 79, 113, 115, 35, 117, 119, 121, 85, 39, 123, 125, 127, 129, 45, 95, 81, 47, 87, 73, 71, 51, 131, 133, 55, 91, 135, 65, 137, 59, 61, 139, 141, 143, 145, 147, 149, 151, 69, 89, 153, 155, 157, 159, 161, 163, 99, 77, 165, 167, 169, 171, 173, 83, 175, 177, 179, 181, 183, 185, 187, 189, 191, 93, 193, 195, 101, 97, 197, 199, 201, 203, 103, 205, 207, 209, 211, 213, 215, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 237, 239, 241, 243, 245, 247, 249, 251, 253, 255, 257, 259, 261, 263, 265, 267, 269, 271, 273, 275, 277, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 341, 343, 345, 347, 349, 351, 353, 355, 357, 359, 361, 363, 365, 367, 369, 371, 373, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 415, 417, 419, 421, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 423, 425, 427, 429, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 431, 433, 435, 437, 439, 441, 443, 445, 447, 449, 451, 453, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 455, 457, 459, 461, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 463, 465, 467, 469, -1, -1, -1, -1, -1, -1, -1, -1, 471, 473, 475, 477, 479, 481, 483, 485, -1, -1, -1, -1, -1, -1, -1, -1, 487, 489, 491, 493, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 10, 6, 8, 16, 22, 36, 14, 12, 122, 98, 20, 30, 24, 18, 34, 38, 62, 50, 72, 102, 26, 52, 28, 76, 120, 86, 54, 32, 46, 56, 92, 114, 44, 124, 40, 42, 100, 48, 180, 134, 194, 90, 130, 60, 224, 156, 132, 68, 64, 174, 58, 96, 66, 88, 110, 70, 198, 226, 82, 162, 78, 168, 74, -1, -1, 94, 190, -1, -1, 80, 228, 188, 144, 128, 152, 146, 216, 84, 230, -1, -1, 212, 210, 126, 196, -1, -1, 106, 206, 232, 104, 136, 118, -1, -1, 234, 142, 236, 116, 108, 238, -1, -1, -1, -1, 240, 112, -1, -1, 242, 244, 148, 246, -1, -1, -1, -1, 178, 248, 250, 158, 140, 252, -1, -1, 166, 172, 214, 164, 222, 138, -1, -1, -1, -1, -1, -1, 218, 160, 154, 254, -1, -1, -1, -1, 256, 150, -1, -1, 184, 258, 260, 262, 186, 264, 266, 268, 270, 200, 176, 272, -1, -1, -1, -1, 170, 274, -1, -1, -1, -1, 204, 276, -1, -1, 202, 278, 182, 280, 282, 208, -1, -1, -1, -1, -1, -1, 284, 192, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 286, 220, -1, -1, -1, -1, 288, 290, -1, -1, 292, 294, 296, 298, -1, -1, 300, 302, -1, -1, 304, 306, 308, 310, -1, -1, -1, -1, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, -1, -1, -1, -1, 332, 334, 336, 338, -1, -1, 340, 342, 344, 346, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 348, 350, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 352, 354, 356, 358, -1, -1, -1, -1, 360, 362, 364, 366, 368, 370, 372, 374, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, -1, -1, -1, -1, -1, -1, -1, -1, 400, 402, 404, 406, 408, 410, 412, 414, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 416, 418, 420, 422, 424, 426, 428, 430, -1, -1, -1, -1, -1, -1, -1, -1, 432, 434, 436, 438, 440, 442, 444, 446, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 12, 18, 48, 10, 54, 26, 16, 22, 14, 36, 30, 60, 70, 20, 40, 138, 212, 24, 106, 72, 34, 200, 28, 52, 96, 32, 64, 80, 232, 44, 90, 206, 38, 112, 104, 120, 42, 188, 100, 46, 328, -1, -1, 50, 184, 148, 94, 178, 144, 56, 290, 158, 58, 216, 128, 134, 62, 76, 142, 152, 66, 68, 88, -1, -1, 78, 298, 194, 74, 86, 166, 84, 172, 156, 116, 308, 82, -1, -1, -1, -1, -1, -1, -1, -1, 92, 224, -1, -1, 236, 244, 98, 252, 182, 170, 330, 102, -1, -1, 114, 234, 256, 108, 110, 124, 118, 332, 162, 334, -1, -1, 268, 336, -1, -1, 174, 122, 146, 164, 126, 316, -1, -1, 130, 338, 132, 340, -1, -1, 136, 228, 168, 250, 302, 140, 342, 344, 226, 346, 198, 348, -1, -1, 350, 150, 352, 354, 154, 262, -1, -1, 222, 248, 280, 160, 240, 356, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 176, 314, -1, -1, 270, 180, -1, -1, -1, -1, 186, 276, 264, 192, 358, 190, -1, -1, 242, 360, 306, 196, -1, -1, -1, -1, 362, 202, 204, 364, 246, 366, 368, 208, 210, 370, -1, -1, 214, 372, 374, 376, 218, 286, 220, 378, -1, -1, -1, -1, -1, -1, -1, -1, 230, 274, -1, -1, 380, 272, -1, -1, 382, 238, -1, -1, 384, 386, -1, -1, 388, 390, -1, -1, -1, -1, -1, -1, 254, 392, -1, -1, 310, 258, 260, 394, -1, -1, -1, -1, 396, 266, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 318, 278, 398, 400, 402, 282, 284, 404, -1, -1, 288, 406, -1, -1, 292, 324, 408, 294, 296, 410, 412, 414, 300, 416, 418, 420, 422, 304, -1, -1, -1, -1, -1, -1, 312, 322, -1, -1, -1, -1, -1, -1, 424, 320, -1, -1, -1, -1, 426, 326, 428, 430, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 432, 434, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 436, 438, -1, -1, -1, -1, 440, 442, -1, -1, -1, -1, 444, 446, 448, 450, -1, -1, 452, 454, -1, -1, 456, 458, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 460, 462, -1, -1, -1, -1, 464, 466, 468, 470, -1, -1, -1, -1, 472, 474, -1, -1, -1, -1, -1, -1, -1, -1, 476, 478, 480, 482, 484, 486, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 488, 490, 492, 494, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 496, 498, 500, 502, -1, -1, -1, -1, -1, -1, -1, -1, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 12, 6, 8, 28, 54, 22, 10, 38, 18, 14, 44, 58, 16, 68, 34, 42, 20, 106, 108, 24, 76, 32, 26, 110, 112, 30, 50, 64, 80, 114, 116, 36, 118, 120, 122, 86, 40, 124, 126, 128, 130, 46, 96, 82, 48, 88, 74, 72, 52, 132, 134, 56, 92, 136, 66, 138, 60, 62, 140, 142, 144, 146, 148, 150, 152, 70, 90, 154, 156, 158, 160, 162, 164, 100, 78, 166, 168, 170, 172, 174, 84, 176, 178, 180, 182, 184, 186, 188, 190, 192, 94, 194, 196, 102, 98, 198, 200, 202, 204, 104, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 424, 426, 428, 430, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 432, 434, 436, 438, 440, 442, 444, 446, 448, 450, 452, 454, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 456, 458, 460, 462, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 464, 466, 468, 470, -1, -1, -1, -1, -1, -1, -1, -1, 472, 474, 476, 478, 480, 482, 484, 486, -1, -1, -1, -1, -1, -1, -1, -1, 488, 490, 492, 494, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 8, 8, 5, 5, 15, 15, 12, 12, 6, 6, 14, 14, 22, 22, 24, 24, 13, 13, 29, 29, 16, 16, 7, 7, 17, 17, 36, 36, 37, 37, 34, 34, 30, 30, 39, 39, 19, 19, 23, 23, 28, 28, 31, 31, 52, 52, 45, 45, 18, 18, 50, 50, 54, 54, 49, 49, 57, 57, 20, 20, 64, 64, 25, 25, 62, 62, 71, 71, 60, 60, 79, 79, 27, 27, 55, 55, 43, 43, 32, 32, 67, 67, 53, 53, 11, 11, 38, 38, 21, 21, 92, 92, 89, 89, 101, 101, 56, 56, 108, 108, 33, 33, 100, 100, 94, 94, 26, 26, 10, 10, 35, 35, 85, 85, 75, 75, 44, 44, 48, 48, 41, 41, 93, 93, 132, 132, 123, 123, 98, 98, 74, 74, 77, 77, 113, 113, 148, 148, 76, 76, 141, 141, 47, 47, 122, 122, 140, 140, 61, 61, 130, 130, 127, 127, 63, 63, 167, 167, 128, 128, 51, 51, 161, 161, 119, 119, 40, 40, 179, 179, 151, 151, 155, 155, 73, 73, 68, 68, 190, 190, 42, 42, 86, 86, 58, 58, 160, 160, 177, 177, 173, 173, 90, 90, 182, 182, 84, 84, 83, 83, 129, 129, 78, 78, 139, 139, 218, 218, 131, 131, 46, 46, 59, 59, 72, 72, 80, 80, 91, 91, 97, 97, 99, 99, 102, 102, 107, 107, 111, 111, 112, 112, 114, 114, 120, 120, 121, 121, 124, 124, 142, 142, 147, 147, 152, 152, 153, 153, 154, 154, 156, 156, 157, 157, 158, 158, 159, 159, 162, 162, 168, 168, 174, 174, 178, 178, 180, 180, 181, 181, 189, 189, 217, 217, 223, 223, 224, 224, 227, 227, 228, 228, 229, 229, 230, 230, 233, 233, 234, 234, 237, 237, 238, 238, 239, 239, 240, 240, 245, 245, 246, 246, 247, 247, 248, 248, 249, 249, 250, 250, 251, 251, 252, 252, 253, 253, 254, 254, 259, 259, 260, 260, 261, 261, 262, 262, 265, 265, 266, 266, 267, 267, 268, 268, 279, 279, 280, 280, 291, 291, 292, 292, 293, 293, 294, 294, 299, 299, 300, 300, 301, 301, 302, 302, 303, 303, 304, 304, 305, 305, 306, 306, 319, 319, 320, 320, 321, 321, 322, 322, 323, 323, 324, 324, 325, 325, 326, 326, 327, 327, 328, 328, 329, 329, 330, 330, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 345, 345, 346, 346, 359, 359, 360, 360, 361, 361, 362, 362, 363, 363, 364, 364, 365, 365, 366, 366, 375, 375, 376, 376, 377, 377, 378, 378, 379, 379, 380, 380, 381, 381, 382, 382, 399, 399, 400, 400, 401, 401, 402, 402, 403, 403, 404, 404, 405, 405, 406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 412, 412, 413, 413, 414, 414, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 4, 4, 12, 12, 10, 10, 5, 5, 17, 17, 11, 11, 21, 21, 9, 9, 26, 26, 14, 14, 29, 29, 24, 24, 13, 13, 36, 36, 18, 18, 40, 40, 33, 33, 43, 43, 6, 6, 47, 47, 27, 27, 8, 8, 53, 53, 56, 56, 15, 15, 60, 60, 30, 30, 64, 64, 65, 65, 16, 16, 23, 23, 72, 72, 61, 61, 69, 69, 31, 31, 80, 80, 75, 75, 73, 73, 66, 66, 34, 34, 89, 89, 50, 50, 28, 28, 95, 95, 42, 42, 100, 100, 38, 38, 22, 22, 106, 106, 107, 107, 37, 37, 103, 103, 78, 78, 109, 109, 39, 39, 120, 120, 108, 108, 123, 123, 58, 58, 127, 127, 129, 129, 59, 59, 133, 133, 19, 19, 138, 138, 62, 62, 52, 52, 121, 121, 49, 49, 148, 148, 63, 63, 151, 151, 77, 77, 55, 55, 158, 158, 111, 111, 122, 122, 74, 74, 135, 135, 98, 98, 76, 76, 119, 119, 173, 173, 51, 51, 178, 178, 97, 97, 48, 48, 183, 183, 41, 41, 188, 188, 186, 186, 71, 71, 194, 194, 143, 143, 25, 25, 200, 200, 201, 201, 35, 35, 206, 206, 207, 207, 20, 20, 211, 211, 57, 57, 215, 215, 217, 217, 155, 155, 90, 90, 141, 141, 134, 134, 227, 227, 32, 32, 104, 104, 93, 93, 236, 236, 159, 159, 191, 191, 94, 94, 203, 203, 156, 156, 136, 136, 96, 96, 251, 251, 105, 105, 256, 256, 257, 257, 152, 152, 185, 185, 264, 264, 115, 115, 177, 177, 232, 232, 228, 228, 184, 184, 276, 276, 157, 157, 280, 280, 281, 281, 216, 216, 285, 285, 54, 54, 289, 289, 292, 292, 293, 293, 70, 70, 297, 297, 137, 137, 302, 302, 193, 193, 79, 79, 255, 255, 309, 309, 174, 174, 124, 124, 275, 275, 318, 318, 310, 310, 290, 290, 324, 324, 44, 44, 99, 99, 110, 110, 112, 112, 116, 116, 128, 128, 130, 130, 139, 139, 140, 140, 142, 142, 144, 144, 147, 147, 149, 149, 150, 150, 160, 160, 187, 187, 192, 192, 199, 199, 202, 202, 204, 204, 205, 205, 208, 208, 212, 212, 213, 213, 214, 214, 218, 218, 231, 231, 235, 235, 239, 239, 240, 240, 243, 243, 244, 244, 252, 252, 258, 258, 263, 263, 277, 277, 278, 278, 279, 279, 282, 282, 286, 286, 291, 291, 294, 294, 295, 295, 296, 296, 298, 298, 299, 299, 300, 300, 301, 301, 317, 317, 323, 323, 325, 325, 326, 326, 337, 337, 338, 338, 349, 349, 350, 350, 355, 355, 356, 356, 361, 361, 362, 362, 363, 363, 364, 364, 367, 367, 368, 368, 371, 371, 372, 372, 401, 401, 402, 402, 407, 407, 408, 408, 409, 409, 410, 410, 415, 415, 416, 416, 425, 425, 426, 426, 427, 427, 428, 428, 429, 429, 430, 430, 443, 443, 444, 444, 445, 445, 446, 446, 463, 463, 464, 464, 465, 465, 466, 466, 475, 475, 476, 476, 477, 477, 478, 478),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 8, 8, 2, 2, 11, 11, 14, 14, 10, 10, 18, 18, 7, 7, 21, 21, 24, 24, 5, 5, 27, 27, 23, 23, 16, 16, 33, 33, 9, 9, 38, 38, 17, 17, 12, 12, 43, 43, 46, 46, 28, 28, 50, 50, 6, 6, 53, 53, 13, 13, 58, 58, 59, 59, 29, 29, 56, 56, 15, 15, 67, 67, 49, 49, 48, 48, 22, 22, 76, 76, 30, 30, 45, 45, 82, 82, 37, 37, 47, 47, 68, 68, 54, 54, 92, 92, 44, 44, 96, 96, 75, 75, 95, 95, 101, 101, 19, 19, 20, 20, 25, 25, 26, 26, 31, 31, 32, 32, 34, 34, 35, 35, 36, 36, 39, 39, 40, 40, 41, 41, 42, 42, 51, 51, 52, 52, 55, 55, 57, 57, 60, 60, 61, 61, 62, 62, 63, 63, 64, 64, 65, 65, 66, 66, 69, 69, 70, 70, 71, 71, 72, 72, 73, 73, 74, 74, 77, 77, 78, 78, 79, 79, 80, 80, 81, 81, 83, 83, 84, 84, 85, 85, 86, 86, 87, 87, 88, 88, 89, 89, 90, 90, 91, 91, 93, 93, 94, 94, 97, 97, 98, 98, 99, 99, 100, 100, 102, 102, 103, 103, 104, 104, 105, 105, 106, 106, 107, 107, 108, 108, 109, 109, 110, 110, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 117, 117, 118, 118, 119, 119, 120, 120, 121, 121, 122, 122, 123, 123, 124, 124, 125, 125, 126, 126, 127, 127, 128, 128, 129, 129, 130, 130, 131, 131, 132, 132, 133, 133, 134, 134, 135, 135, 136, 136, 137, 137, 138, 138, 139, 139, 140, 140, 141, 141, 142, 142, 143, 143, 144, 144, 145, 145, 146, 146, 147, 147, 148, 148, 149, 149, 150, 150, 151, 151, 152, 152, 153, 153, 154, 154, 155, 155, 156, 156, 157, 157, 158, 158, 159, 159, 160, 160, 161, 161, 162, 162, 163, 163, 164, 164, 165, 165, 166, 166, 167, 167, 168, 168, 169, 169, 170, 170, 171, 171, 172, 172, 173, 173, 174, 174, 175, 175, 176, 176, 177, 177, 178, 178, 179, 179, 180, 180, 181, 181, 182, 182, 183, 183, 184, 184, 185, 185, 186, 186, 187, 187, 188, 188, 189, 189, 190, 190, 191, 191, 192, 192, 193, 193, 194, 194, 195, 195, 196, 196, 197, 197, 198, 198, 199, 199, 200, 200, 201, 201, 202, 202, 203, 203, 204, 204, 205, 205, 206, 206, 207, 207, 208, 208, 209, 209, 210, 210, 235, 235, 236, 236, 237, 237, 238, 238, 271, 271, 272, 272, 273, 273, 274, 274, 275, 275, 276, 276, 277, 277, 278, 278, 279, 279, 280, 280, 281, 281, 282, 282, 347, 347, 348, 348, 349, 349, 350, 350, 383, 383, 384, 384, 385, 385, 386, 386, 395, 395, 396, 396, 397, 397, 398, 398, 399, 399, 400, 400, 401, 401, 402, 402, 411, 411, 412, 412, 413, 413, 414, 414, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 5, 5, 6, 6, 5, 5, 4, 4, 6, 6, 5, 5, 7, 7, 6, 6, 6, 6, 6, 6, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 8, 8, 6, 6, 8, 8, 5, 5, 7, 7, 6, 6, 7, 7, 6, 6, 8, 8, 7, 7, 7, 7, 8, 8, 7, 7, 7, 7, 7, 7, 8, 8, 4, 4, 7, 7, 5, 5, 8, 8, 8, 8, 6, 6, 8, 8, 7, 7, 6, 6, 8, 8, 8, 8, 6, 6, 3, 3, 5, 5, 8, 8, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 6, 6, 5, 5, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 6, 6, 7, 7, 4, 4, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 5, 5, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 4, 4, 6, 6, 6, 6, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 5, 5, 5, 5, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 5, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 6, 6, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 6, 6, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 5, 5, 6, 6, 5, 5, 6, 6, 7, 7, 8, 8, 4, 4, 5, 5, 6, 6, 3, 3, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 5, 5, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 4, 4, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 5, 5, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 4, 4, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6, 4, 4, 5, 5, 6, 6, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 5, 5, 6, 6, 6, 6, 3, 3, 4, 4, 5, 5, 5, 5, 6, 6, 4, 4, 5, 5, 4, 4, 5, 5, 6, 6, 6, 6, 6, 6, 5, 5, 6, 6, 6, 6, 6, 6, 5, 5, 6, 6, 6, 6, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 5, 5, 6, 6, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 6, 6, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((65, 66, 69, 70, 81, 82, 87, 88, 95, 96, 103, 104, 105, 106, 109, 110, 115, 116, 117, 118, 125, 126, 133, 134, 135, 136, 137, 138, 143, 144, 145, 146, 149, 150, 163, 164, 165, 166, 169, 170, 171, 172, 175, 176, 183, 184, 185, 186, 187, 188, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 219, 220, 221, 222, 225, 226, 231, 232, 235, 236, 241, 242, 243, 244, 255, 256, 257, 258, 263, 264, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 295, 296, 297, 298, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 331, 332, 333, 334, 335, 336, 337, 338, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 367, 368, 369, 370, 371, 372, 373, 374, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510),
                (45, 46, 67, 68, 81, 82, 83, 84, 85, 86, 87, 88, 91, 92, 101, 102, 113, 114, 117, 118, 125, 126, 131, 132, 145, 146, 153, 154, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 175, 176, 179, 180, 181, 182, 189, 190, 195, 196, 197, 198, 209, 210, 219, 220, 221, 222, 223, 224, 225, 226, 229, 230, 233, 234, 237, 238, 241, 242, 245, 246, 247, 248, 249, 250, 253, 254, 259, 260, 261, 262, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 283, 284, 287, 288, 303, 304, 305, 306, 307, 308, 311, 312, 313, 314, 315, 316, 319, 320, 321, 322, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 351, 352, 353, 354, 357, 358, 359, 360, 365, 366, 369, 370, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 403, 404, 405, 406, 411, 412, 413, 414, 417, 418, 419, 420, 421, 422, 423, 424, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 467, 468, 469, 470, 471, 472, 473, 474, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510),
                (211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 387, 388, 389, 390, 391, 392, 393, 394, 403, 404, 405, 406, 407, 408, 409, 410, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
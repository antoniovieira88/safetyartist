library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 2, 0, 0, -2, -2, 2, -2, -2, 1, 2, -2, -2, 2, -2, -2, 1, 1, 2, -2, -2, 1, -2, -2, 1, 2, -2, -2, 2, -2, -2),
                (0, 2, 0, 1, -2, -2, 0, -2, -2, 0, 0, -2, -2, 2, -2, -2, 1, 1, 1, -2, -2, 0, -2, -2, 2, 2, -2, -2, 1, -2, -2),
                (1, 1, 2, 0, -2, -2, 1, -2, -2, 1, 0, -2, -2, 2, -2, -2, 0, 0, 1, -2, -2, 0, -2, -2, 0, 2, -2, -2, 0, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((34460, 134, 16405, 3670, -256, -256, 109, -256, -256, 1771, 164, -256, -256, 164, -256, -256, 3039, 2709, 92, -256, -256, 2709, -256, -256, 3395, 134, -256, -256, 134, -256, -256),
                (34460, 134, 12612, 920, -256, -256, 24386, -256, -256, 10276, 6389, -256, -256, 164, -256, -256, 3029, 2693, 2419, -256, -256, 47292, -256, -256, 134, 109, -256, -256, 3518, -256, -256),
                (2202, 1444, 109, 10323, -256, -256, 827, -256, -256, 1773, 17571, -256, -256, 92, -256, -256, 44659, 34513, 2580, -256, -256, 39576, -256, -256, 66386, 109, -256, -256, 77116, -256, -256)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((38, 18, 17, 10, 3, 13, 23, 22, 25, 20, 34, 34, 35, 7, 6, 7, 42, 42, 43, 42, 43, 41, 0, 41, 38, 38, 37, 41, 36, 35, 39),
                (38, 18, 17, 8, 29, 1, 22, 19, 25, 20, 9, 5, 14, 25, 24, 27, 42, 42, 43, 43, 42, 41, 18, 42, 38, 36, 35, 38, 40, 41, 38),
                (38, 41, 42, 41, 17, 43, 42, 42, 41, 39, 40, 3, 42, 38, 37, 39, 35, 4, 1, 3, 0, 16, 13, 18, 41, 30, 21, 37, 42, 38, 43)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
-------------------------------------------------------------------
-- File   : rom_4096x16.vhd
-------------------------------------------------------------------
-- Descricao : Synchronous 4096x16 ROM.
-------------------------------------------------------------------
-- Revision:
--     Date        Rev     Author            Description
--     05/07/2023  1.0     Antonio V.S.Neto  Creation.
-------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_4096x16 is
   port (
       address   : in  std_logic_vector(11 downto 0);
	   clk       : in  std_logic;
       out_rom   : out std_logic_vector(15 downto 0)
    );
end entity rom_4096x16;

-- Initial data explicitly declared 
architecture rom_bcd of rom_4096x16 is
  type   memory_struct is array(0 to 4095) of std_logic_vector(15 downto 0);
  signal memory : memory_struct := (
									"0000000000000000",
									"0000000000000001",
									"0000000000000010",
									"0000000000000011",
									"0000000000000100",
									"0000000000000101",
									"0000000000000110",
									"0000000000000111",
									"0000000000001000",
									"0000000000001001",
									"0000000000010000",
									"0000000000010001",
									"0000000000010010",
									"0000000000010011",
									"0000000000010100",
									"0000000000010101",
									"0000000000010110",
									"0000000000010111",
									"0000000000011000",
									"0000000000011001",
									"0000000000100000",
									"0000000000100001",
									"0000000000100010",
									"0000000000100011",
									"0000000000100100",
									"0000000000100101",
									"0000000000100110",
									"0000000000100111",
									"0000000000101000",
									"0000000000101001",
									"0000000000110000",
									"0000000000110001",
									"0000000000110010",
									"0000000000110011",
									"0000000000110100",
									"0000000000110101",
									"0000000000110110",
									"0000000000110111",
									"0000000000111000",
									"0000000000111001",
									"0000000001000000",
									"0000000001000001",
									"0000000001000010",
									"0000000001000011",
									"0000000001000100",
									"0000000001000101",
									"0000000001000110",
									"0000000001000111",
									"0000000001001000",
									"0000000001001001",
									"0000000001010000",
									"0000000001010001",
									"0000000001010010",
									"0000000001010011",
									"0000000001010100",
									"0000000001010101",
									"0000000001010110",
									"0000000001010111",
									"0000000001011000",
									"0000000001011001",
									"0000000001100000",
									"0000000001100001",
									"0000000001100010",
									"0000000001100011",
									"0000000001100100",
									"0000000001100101",
									"0000000001100110",
									"0000000001100111",
									"0000000001101000",
									"0000000001101001",
									"0000000001110000",
									"0000000001110001",
									"0000000001110010",
									"0000000001110011",
									"0000000001110100",
									"0000000001110101",
									"0000000001110110",
									"0000000001110111",
									"0000000001111000",
									"0000000001111001",
									"0000000010000000",
									"0000000010000001",
									"0000000010000010",
									"0000000010000011",
									"0000000010000100",
									"0000000010000101",
									"0000000010000110",
									"0000000010000111",
									"0000000010001000",
									"0000000010001001",
									"0000000010010000",
									"0000000010010001",
									"0000000010010010",
									"0000000010010011",
									"0000000010010100",
									"0000000010010101",
									"0000000010010110",
									"0000000010010111",
									"0000000010011000",
									"0000000010011001",
									"0000000100000000",
									"0000000100000001",
									"0000000100000010",
									"0000000100000011",
									"0000000100000100",
									"0000000100000101",
									"0000000100000110",
									"0000000100000111",
									"0000000100001000",
									"0000000100001001",
									"0000000100010000",
									"0000000100010001",
									"0000000100010010",
									"0000000100010011",
									"0000000100010100",
									"0000000100010101",
									"0000000100010110",
									"0000000100010111",
									"0000000100011000",
									"0000000100011001",
									"0000000100100000",
									"0000000100100001",
									"0000000100100010",
									"0000000100100011",
									"0000000100100100",
									"0000000100100101",
									"0000000100100110",
									"0000000100100111",
									"0000000100101000",
									"0000000100101001",
									"0000000100110000",
									"0000000100110001",
									"0000000100110010",
									"0000000100110011",
									"0000000100110100",
									"0000000100110101",
									"0000000100110110",
									"0000000100110111",
									"0000000100111000",
									"0000000100111001",
									"0000000101000000",
									"0000000101000001",
									"0000000101000010",
									"0000000101000011",
									"0000000101000100",
									"0000000101000101",
									"0000000101000110",
									"0000000101000111",
									"0000000101001000",
									"0000000101001001",
									"0000000101010000",
									"0000000101010001",
									"0000000101010010",
									"0000000101010011",
									"0000000101010100",
									"0000000101010101",
									"0000000101010110",
									"0000000101010111",
									"0000000101011000",
									"0000000101011001",
									"0000000101100000",
									"0000000101100001",
									"0000000101100010",
									"0000000101100011",
									"0000000101100100",
									"0000000101100101",
									"0000000101100110",
									"0000000101100111",
									"0000000101101000",
									"0000000101101001",
									"0000000101110000",
									"0000000101110001",
									"0000000101110010",
									"0000000101110011",
									"0000000101110100",
									"0000000101110101",
									"0000000101110110",
									"0000000101110111",
									"0000000101111000",
									"0000000101111001",
									"0000000110000000",
									"0000000110000001",
									"0000000110000010",
									"0000000110000011",
									"0000000110000100",
									"0000000110000101",
									"0000000110000110",
									"0000000110000111",
									"0000000110001000",
									"0000000110001001",
									"0000000110010000",
									"0000000110010001",
									"0000000110010010",
									"0000000110010011",
									"0000000110010100",
									"0000000110010101",
									"0000000110010110",
									"0000000110010111",
									"0000000110011000",
									"0000000110011001",
									"0000001000000000",
									"0000001000000001",
									"0000001000000010",
									"0000001000000011",
									"0000001000000100",
									"0000001000000101",
									"0000001000000110",
									"0000001000000111",
									"0000001000001000",
									"0000001000001001",
									"0000001000010000",
									"0000001000010001",
									"0000001000010010",
									"0000001000010011",
									"0000001000010100",
									"0000001000010101",
									"0000001000010110",
									"0000001000010111",
									"0000001000011000",
									"0000001000011001",
									"0000001000100000",
									"0000001000100001",
									"0000001000100010",
									"0000001000100011",
									"0000001000100100",
									"0000001000100101",
									"0000001000100110",
									"0000001000100111",
									"0000001000101000",
									"0000001000101001",
									"0000001000110000",
									"0000001000110001",
									"0000001000110010",
									"0000001000110011",
									"0000001000110100",
									"0000001000110101",
									"0000001000110110",
									"0000001000110111",
									"0000001000111000",
									"0000001000111001",
									"0000001001000000",
									"0000001001000001",
									"0000001001000010",
									"0000001001000011",
									"0000001001000100",
									"0000001001000101",
									"0000001001000110",
									"0000001001000111",
									"0000001001001000",
									"0000001001001001",
									"0000001001010000",
									"0000001001010001",
									"0000001001010010",
									"0000001001010011",
									"0000001001010100",
									"0000001001010101",
									"0000001001010110",
									"0000001001010111",
									"0000001001011000",
									"0000001001011001",
									"0000001001100000",
									"0000001001100001",
									"0000001001100010",
									"0000001001100011",
									"0000001001100100",
									"0000001001100101",
									"0000001001100110",
									"0000001001100111",
									"0000001001101000",
									"0000001001101001",
									"0000001001110000",
									"0000001001110001",
									"0000001001110010",
									"0000001001110011",
									"0000001001110100",
									"0000001001110101",
									"0000001001110110",
									"0000001001110111",
									"0000001001111000",
									"0000001001111001",
									"0000001010000000",
									"0000001010000001",
									"0000001010000010",
									"0000001010000011",
									"0000001010000100",
									"0000001010000101",
									"0000001010000110",
									"0000001010000111",
									"0000001010001000",
									"0000001010001001",
									"0000001010010000",
									"0000001010010001",
									"0000001010010010",
									"0000001010010011",
									"0000001010010100",
									"0000001010010101",
									"0000001010010110",
									"0000001010010111",
									"0000001010011000",
									"0000001010011001",
									"0000001100000000",
									"0000001100000001",
									"0000001100000010",
									"0000001100000011",
									"0000001100000100",
									"0000001100000101",
									"0000001100000110",
									"0000001100000111",
									"0000001100001000",
									"0000001100001001",
									"0000001100010000",
									"0000001100010001",
									"0000001100010010",
									"0000001100010011",
									"0000001100010100",
									"0000001100010101",
									"0000001100010110",
									"0000001100010111",
									"0000001100011000",
									"0000001100011001",
									"0000001100100000",
									"0000001100100001",
									"0000001100100010",
									"0000001100100011",
									"0000001100100100",
									"0000001100100101",
									"0000001100100110",
									"0000001100100111",
									"0000001100101000",
									"0000001100101001",
									"0000001100110000",
									"0000001100110001",
									"0000001100110010",
									"0000001100110011",
									"0000001100110100",
									"0000001100110101",
									"0000001100110110",
									"0000001100110111",
									"0000001100111000",
									"0000001100111001",
									"0000001101000000",
									"0000001101000001",
									"0000001101000010",
									"0000001101000011",
									"0000001101000100",
									"0000001101000101",
									"0000001101000110",
									"0000001101000111",
									"0000001101001000",
									"0000001101001001",
									"0000001101010000",
									"0000001101010001",
									"0000001101010010",
									"0000001101010011",
									"0000001101010100",
									"0000001101010101",
									"0000001101010110",
									"0000001101010111",
									"0000001101011000",
									"0000001101011001",
									"0000001101100000",
									"0000001101100001",
									"0000001101100010",
									"0000001101100011",
									"0000001101100100",
									"0000001101100101",
									"0000001101100110",
									"0000001101100111",
									"0000001101101000",
									"0000001101101001",
									"0000001101110000",
									"0000001101110001",
									"0000001101110010",
									"0000001101110011",
									"0000001101110100",
									"0000001101110101",
									"0000001101110110",
									"0000001101110111",
									"0000001101111000",
									"0000001101111001",
									"0000001110000000",
									"0000001110000001",
									"0000001110000010",
									"0000001110000011",
									"0000001110000100",
									"0000001110000101",
									"0000001110000110",
									"0000001110000111",
									"0000001110001000",
									"0000001110001001",
									"0000001110010000",
									"0000001110010001",
									"0000001110010010",
									"0000001110010011",
									"0000001110010100",
									"0000001110010101",
									"0000001110010110",
									"0000001110010111",
									"0000001110011000",
									"0000001110011001",
									"0000010000000000",
									"0000010000000001",
									"0000010000000010",
									"0000010000000011",
									"0000010000000100",
									"0000010000000101",
									"0000010000000110",
									"0000010000000111",
									"0000010000001000",
									"0000010000001001",
									"0000010000010000",
									"0000010000010001",
									"0000010000010010",
									"0000010000010011",
									"0000010000010100",
									"0000010000010101",
									"0000010000010110",
									"0000010000010111",
									"0000010000011000",
									"0000010000011001",
									"0000010000100000",
									"0000010000100001",
									"0000010000100010",
									"0000010000100011",
									"0000010000100100",
									"0000010000100101",
									"0000010000100110",
									"0000010000100111",
									"0000010000101000",
									"0000010000101001",
									"0000010000110000",
									"0000010000110001",
									"0000010000110010",
									"0000010000110011",
									"0000010000110100",
									"0000010000110101",
									"0000010000110110",
									"0000010000110111",
									"0000010000111000",
									"0000010000111001",
									"0000010001000000",
									"0000010001000001",
									"0000010001000010",
									"0000010001000011",
									"0000010001000100",
									"0000010001000101",
									"0000010001000110",
									"0000010001000111",
									"0000010001001000",
									"0000010001001001",
									"0000010001010000",
									"0000010001010001",
									"0000010001010010",
									"0000010001010011",
									"0000010001010100",
									"0000010001010101",
									"0000010001010110",
									"0000010001010111",
									"0000010001011000",
									"0000010001011001",
									"0000010001100000",
									"0000010001100001",
									"0000010001100010",
									"0000010001100011",
									"0000010001100100",
									"0000010001100101",
									"0000010001100110",
									"0000010001100111",
									"0000010001101000",
									"0000010001101001",
									"0000010001110000",
									"0000010001110001",
									"0000010001110010",
									"0000010001110011",
									"0000010001110100",
									"0000010001110101",
									"0000010001110110",
									"0000010001110111",
									"0000010001111000",
									"0000010001111001",
									"0000010010000000",
									"0000010010000001",
									"0000010010000010",
									"0000010010000011",
									"0000010010000100",
									"0000010010000101",
									"0000010010000110",
									"0000010010000111",
									"0000010010001000",
									"0000010010001001",
									"0000010010010000",
									"0000010010010001",
									"0000010010010010",
									"0000010010010011",
									"0000010010010100",
									"0000010010010101",
									"0000010010010110",
									"0000010010010111",
									"0000010010011000",
									"0000010010011001",
									"0000010100000000",
									"0000010100000001",
									"0000010100000010",
									"0000010100000011",
									"0000010100000100",
									"0000010100000101",
									"0000010100000110",
									"0000010100000111",
									"0000010100001000",
									"0000010100001001",
									"0000010100010000",
									"0000010100010001",
									"0000010100010010",
									"0000010100010011",
									"0000010100010100",
									"0000010100010101",
									"0000010100010110",
									"0000010100010111",
									"0000010100011000",
									"0000010100011001",
									"0000010100100000",
									"0000010100100001",
									"0000010100100010",
									"0000010100100011",
									"0000010100100100",
									"0000010100100101",
									"0000010100100110",
									"0000010100100111",
									"0000010100101000",
									"0000010100101001",
									"0000010100110000",
									"0000010100110001",
									"0000010100110010",
									"0000010100110011",
									"0000010100110100",
									"0000010100110101",
									"0000010100110110",
									"0000010100110111",
									"0000010100111000",
									"0000010100111001",
									"0000010101000000",
									"0000010101000001",
									"0000010101000010",
									"0000010101000011",
									"0000010101000100",
									"0000010101000101",
									"0000010101000110",
									"0000010101000111",
									"0000010101001000",
									"0000010101001001",
									"0000010101010000",
									"0000010101010001",
									"0000010101010010",
									"0000010101010011",
									"0000010101010100",
									"0000010101010101",
									"0000010101010110",
									"0000010101010111",
									"0000010101011000",
									"0000010101011001",
									"0000010101100000",
									"0000010101100001",
									"0000010101100010",
									"0000010101100011",
									"0000010101100100",
									"0000010101100101",
									"0000010101100110",
									"0000010101100111",
									"0000010101101000",
									"0000010101101001",
									"0000010101110000",
									"0000010101110001",
									"0000010101110010",
									"0000010101110011",
									"0000010101110100",
									"0000010101110101",
									"0000010101110110",
									"0000010101110111",
									"0000010101111000",
									"0000010101111001",
									"0000010110000000",
									"0000010110000001",
									"0000010110000010",
									"0000010110000011",
									"0000010110000100",
									"0000010110000101",
									"0000010110000110",
									"0000010110000111",
									"0000010110001000",
									"0000010110001001",
									"0000010110010000",
									"0000010110010001",
									"0000010110010010",
									"0000010110010011",
									"0000010110010100",
									"0000010110010101",
									"0000010110010110",
									"0000010110010111",
									"0000010110011000",
									"0000010110011001",
									"0000011000000000",
									"0000011000000001",
									"0000011000000010",
									"0000011000000011",
									"0000011000000100",
									"0000011000000101",
									"0000011000000110",
									"0000011000000111",
									"0000011000001000",
									"0000011000001001",
									"0000011000010000",
									"0000011000010001",
									"0000011000010010",
									"0000011000010011",
									"0000011000010100",
									"0000011000010101",
									"0000011000010110",
									"0000011000010111",
									"0000011000011000",
									"0000011000011001",
									"0000011000100000",
									"0000011000100001",
									"0000011000100010",
									"0000011000100011",
									"0000011000100100",
									"0000011000100101",
									"0000011000100110",
									"0000011000100111",
									"0000011000101000",
									"0000011000101001",
									"0000011000110000",
									"0000011000110001",
									"0000011000110010",
									"0000011000110011",
									"0000011000110100",
									"0000011000110101",
									"0000011000110110",
									"0000011000110111",
									"0000011000111000",
									"0000011000111001",
									"0000011001000000",
									"0000011001000001",
									"0000011001000010",
									"0000011001000011",
									"0000011001000100",
									"0000011001000101",
									"0000011001000110",
									"0000011001000111",
									"0000011001001000",
									"0000011001001001",
									"0000011001010000",
									"0000011001010001",
									"0000011001010010",
									"0000011001010011",
									"0000011001010100",
									"0000011001010101",
									"0000011001010110",
									"0000011001010111",
									"0000011001011000",
									"0000011001011001",
									"0000011001100000",
									"0000011001100001",
									"0000011001100010",
									"0000011001100011",
									"0000011001100100",
									"0000011001100101",
									"0000011001100110",
									"0000011001100111",
									"0000011001101000",
									"0000011001101001",
									"0000011001110000",
									"0000011001110001",
									"0000011001110010",
									"0000011001110011",
									"0000011001110100",
									"0000011001110101",
									"0000011001110110",
									"0000011001110111",
									"0000011001111000",
									"0000011001111001",
									"0000011010000000",
									"0000011010000001",
									"0000011010000010",
									"0000011010000011",
									"0000011010000100",
									"0000011010000101",
									"0000011010000110",
									"0000011010000111",
									"0000011010001000",
									"0000011010001001",
									"0000011010010000",
									"0000011010010001",
									"0000011010010010",
									"0000011010010011",
									"0000011010010100",
									"0000011010010101",
									"0000011010010110",
									"0000011010010111",
									"0000011010011000",
									"0000011010011001",
									"0000011100000000",
									"0000011100000001",
									"0000011100000010",
									"0000011100000011",
									"0000011100000100",
									"0000011100000101",
									"0000011100000110",
									"0000011100000111",
									"0000011100001000",
									"0000011100001001",
									"0000011100010000",
									"0000011100010001",
									"0000011100010010",
									"0000011100010011",
									"0000011100010100",
									"0000011100010101",
									"0000011100010110",
									"0000011100010111",
									"0000011100011000",
									"0000011100011001",
									"0000011100100000",
									"0000011100100001",
									"0000011100100010",
									"0000011100100011",
									"0000011100100100",
									"0000011100100101",
									"0000011100100110",
									"0000011100100111",
									"0000011100101000",
									"0000011100101001",
									"0000011100110000",
									"0000011100110001",
									"0000011100110010",
									"0000011100110011",
									"0000011100110100",
									"0000011100110101",
									"0000011100110110",
									"0000011100110111",
									"0000011100111000",
									"0000011100111001",
									"0000011101000000",
									"0000011101000001",
									"0000011101000010",
									"0000011101000011",
									"0000011101000100",
									"0000011101000101",
									"0000011101000110",
									"0000011101000111",
									"0000011101001000",
									"0000011101001001",
									"0000011101010000",
									"0000011101010001",
									"0000011101010010",
									"0000011101010011",
									"0000011101010100",
									"0000011101010101",
									"0000011101010110",
									"0000011101010111",
									"0000011101011000",
									"0000011101011001",
									"0000011101100000",
									"0000011101100001",
									"0000011101100010",
									"0000011101100011",
									"0000011101100100",
									"0000011101100101",
									"0000011101100110",
									"0000011101100111",
									"0000011101101000",
									"0000011101101001",
									"0000011101110000",
									"0000011101110001",
									"0000011101110010",
									"0000011101110011",
									"0000011101110100",
									"0000011101110101",
									"0000011101110110",
									"0000011101110111",
									"0000011101111000",
									"0000011101111001",
									"0000011110000000",
									"0000011110000001",
									"0000011110000010",
									"0000011110000011",
									"0000011110000100",
									"0000011110000101",
									"0000011110000110",
									"0000011110000111",
									"0000011110001000",
									"0000011110001001",
									"0000011110010000",
									"0000011110010001",
									"0000011110010010",
									"0000011110010011",
									"0000011110010100",
									"0000011110010101",
									"0000011110010110",
									"0000011110010111",
									"0000011110011000",
									"0000011110011001",
									"0000100000000000",
									"0000100000000001",
									"0000100000000010",
									"0000100000000011",
									"0000100000000100",
									"0000100000000101",
									"0000100000000110",
									"0000100000000111",
									"0000100000001000",
									"0000100000001001",
									"0000100000010000",
									"0000100000010001",
									"0000100000010010",
									"0000100000010011",
									"0000100000010100",
									"0000100000010101",
									"0000100000010110",
									"0000100000010111",
									"0000100000011000",
									"0000100000011001",
									"0000100000100000",
									"0000100000100001",
									"0000100000100010",
									"0000100000100011",
									"0000100000100100",
									"0000100000100101",
									"0000100000100110",
									"0000100000100111",
									"0000100000101000",
									"0000100000101001",
									"0000100000110000",
									"0000100000110001",
									"0000100000110010",
									"0000100000110011",
									"0000100000110100",
									"0000100000110101",
									"0000100000110110",
									"0000100000110111",
									"0000100000111000",
									"0000100000111001",
									"0000100001000000",
									"0000100001000001",
									"0000100001000010",
									"0000100001000011",
									"0000100001000100",
									"0000100001000101",
									"0000100001000110",
									"0000100001000111",
									"0000100001001000",
									"0000100001001001",
									"0000100001010000",
									"0000100001010001",
									"0000100001010010",
									"0000100001010011",
									"0000100001010100",
									"0000100001010101",
									"0000100001010110",
									"0000100001010111",
									"0000100001011000",
									"0000100001011001",
									"0000100001100000",
									"0000100001100001",
									"0000100001100010",
									"0000100001100011",
									"0000100001100100",
									"0000100001100101",
									"0000100001100110",
									"0000100001100111",
									"0000100001101000",
									"0000100001101001",
									"0000100001110000",
									"0000100001110001",
									"0000100001110010",
									"0000100001110011",
									"0000100001110100",
									"0000100001110101",
									"0000100001110110",
									"0000100001110111",
									"0000100001111000",
									"0000100001111001",
									"0000100010000000",
									"0000100010000001",
									"0000100010000010",
									"0000100010000011",
									"0000100010000100",
									"0000100010000101",
									"0000100010000110",
									"0000100010000111",
									"0000100010001000",
									"0000100010001001",
									"0000100010010000",
									"0000100010010001",
									"0000100010010010",
									"0000100010010011",
									"0000100010010100",
									"0000100010010101",
									"0000100010010110",
									"0000100010010111",
									"0000100010011000",
									"0000100010011001",
									"0000100100000000",
									"0000100100000001",
									"0000100100000010",
									"0000100100000011",
									"0000100100000100",
									"0000100100000101",
									"0000100100000110",
									"0000100100000111",
									"0000100100001000",
									"0000100100001001",
									"0000100100010000",
									"0000100100010001",
									"0000100100010010",
									"0000100100010011",
									"0000100100010100",
									"0000100100010101",
									"0000100100010110",
									"0000100100010111",
									"0000100100011000",
									"0000100100011001",
									"0000100100100000",
									"0000100100100001",
									"0000100100100010",
									"0000100100100011",
									"0000100100100100",
									"0000100100100101",
									"0000100100100110",
									"0000100100100111",
									"0000100100101000",
									"0000100100101001",
									"0000100100110000",
									"0000100100110001",
									"0000100100110010",
									"0000100100110011",
									"0000100100110100",
									"0000100100110101",
									"0000100100110110",
									"0000100100110111",
									"0000100100111000",
									"0000100100111001",
									"0000100101000000",
									"0000100101000001",
									"0000100101000010",
									"0000100101000011",
									"0000100101000100",
									"0000100101000101",
									"0000100101000110",
									"0000100101000111",
									"0000100101001000",
									"0000100101001001",
									"0000100101010000",
									"0000100101010001",
									"0000100101010010",
									"0000100101010011",
									"0000100101010100",
									"0000100101010101",
									"0000100101010110",
									"0000100101010111",
									"0000100101011000",
									"0000100101011001",
									"0000100101100000",
									"0000100101100001",
									"0000100101100010",
									"0000100101100011",
									"0000100101100100",
									"0000100101100101",
									"0000100101100110",
									"0000100101100111",
									"0000100101101000",
									"0000100101101001",
									"0000100101110000",
									"0000100101110001",
									"0000100101110010",
									"0000100101110011",
									"0000100101110100",
									"0000100101110101",
									"0000100101110110",
									"0000100101110111",
									"0000100101111000",
									"0000100101111001",
									"0000100110000000",
									"0000100110000001",
									"0000100110000010",
									"0000100110000011",
									"0000100110000100",
									"0000100110000101",
									"0000100110000110",
									"0000100110000111",
									"0000100110001000",
									"0000100110001001",
									"0000100110010000",
									"0000100110010001",
									"0000100110010010",
									"0000100110010011",
									"0000100110010100",
									"0000100110010101",
									"0000100110010110",
									"0000100110010111",
									"0000100110011000",
									"0000100110011001",
									"0001000000000000",
									"0001000000000001",
									"0001000000000010",
									"0001000000000011",
									"0001000000000100",
									"0001000000000101",
									"0001000000000110",
									"0001000000000111",
									"0001000000001000",
									"0001000000001001",
									"0001000000010000",
									"0001000000010001",
									"0001000000010010",
									"0001000000010011",
									"0001000000010100",
									"0001000000010101",
									"0001000000010110",
									"0001000000010111",
									"0001000000011000",
									"0001000000011001",
									"0001000000100000",
									"0001000000100001",
									"0001000000100010",
									"0001000000100011",
									"0001000000100100",
									"0001000000100101",
									"0001000000100110",
									"0001000000100111",
									"0001000000101000",
									"0001000000101001",
									"0001000000110000",
									"0001000000110001",
									"0001000000110010",
									"0001000000110011",
									"0001000000110100",
									"0001000000110101",
									"0001000000110110",
									"0001000000110111",
									"0001000000111000",
									"0001000000111001",
									"0001000001000000",
									"0001000001000001",
									"0001000001000010",
									"0001000001000011",
									"0001000001000100",
									"0001000001000101",
									"0001000001000110",
									"0001000001000111",
									"0001000001001000",
									"0001000001001001",
									"0001000001010000",
									"0001000001010001",
									"0001000001010010",
									"0001000001010011",
									"0001000001010100",
									"0001000001010101",
									"0001000001010110",
									"0001000001010111",
									"0001000001011000",
									"0001000001011001",
									"0001000001100000",
									"0001000001100001",
									"0001000001100010",
									"0001000001100011",
									"0001000001100100",
									"0001000001100101",
									"0001000001100110",
									"0001000001100111",
									"0001000001101000",
									"0001000001101001",
									"0001000001110000",
									"0001000001110001",
									"0001000001110010",
									"0001000001110011",
									"0001000001110100",
									"0001000001110101",
									"0001000001110110",
									"0001000001110111",
									"0001000001111000",
									"0001000001111001",
									"0001000010000000",
									"0001000010000001",
									"0001000010000010",
									"0001000010000011",
									"0001000010000100",
									"0001000010000101",
									"0001000010000110",
									"0001000010000111",
									"0001000010001000",
									"0001000010001001",
									"0001000010010000",
									"0001000010010001",
									"0001000010010010",
									"0001000010010011",
									"0001000010010100",
									"0001000010010101",
									"0001000010010110",
									"0001000010010111",
									"0001000010011000",
									"0001000010011001",
									"0001000100000000",
									"0001000100000001",
									"0001000100000010",
									"0001000100000011",
									"0001000100000100",
									"0001000100000101",
									"0001000100000110",
									"0001000100000111",
									"0001000100001000",
									"0001000100001001",
									"0001000100010000",
									"0001000100010001",
									"0001000100010010",
									"0001000100010011",
									"0001000100010100",
									"0001000100010101",
									"0001000100010110",
									"0001000100010111",
									"0001000100011000",
									"0001000100011001",
									"0001000100100000",
									"0001000100100001",
									"0001000100100010",
									"0001000100100011",
									"0001000100100100",
									"0001000100100101",
									"0001000100100110",
									"0001000100100111",
									"0001000100101000",
									"0001000100101001",
									"0001000100110000",
									"0001000100110001",
									"0001000100110010",
									"0001000100110011",
									"0001000100110100",
									"0001000100110101",
									"0001000100110110",
									"0001000100110111",
									"0001000100111000",
									"0001000100111001",
									"0001000101000000",
									"0001000101000001",
									"0001000101000010",
									"0001000101000011",
									"0001000101000100",
									"0001000101000101",
									"0001000101000110",
									"0001000101000111",
									"0001000101001000",
									"0001000101001001",
									"0001000101010000",
									"0001000101010001",
									"0001000101010010",
									"0001000101010011",
									"0001000101010100",
									"0001000101010101",
									"0001000101010110",
									"0001000101010111",
									"0001000101011000",
									"0001000101011001",
									"0001000101100000",
									"0001000101100001",
									"0001000101100010",
									"0001000101100011",
									"0001000101100100",
									"0001000101100101",
									"0001000101100110",
									"0001000101100111",
									"0001000101101000",
									"0001000101101001",
									"0001000101110000",
									"0001000101110001",
									"0001000101110010",
									"0001000101110011",
									"0001000101110100",
									"0001000101110101",
									"0001000101110110",
									"0001000101110111",
									"0001000101111000",
									"0001000101111001",
									"0001000110000000",
									"0001000110000001",
									"0001000110000010",
									"0001000110000011",
									"0001000110000100",
									"0001000110000101",
									"0001000110000110",
									"0001000110000111",
									"0001000110001000",
									"0001000110001001",
									"0001000110010000",
									"0001000110010001",
									"0001000110010010",
									"0001000110010011",
									"0001000110010100",
									"0001000110010101",
									"0001000110010110",
									"0001000110010111",
									"0001000110011000",
									"0001000110011001",
									"0001001000000000",
									"0001001000000001",
									"0001001000000010",
									"0001001000000011",
									"0001001000000100",
									"0001001000000101",
									"0001001000000110",
									"0001001000000111",
									"0001001000001000",
									"0001001000001001",
									"0001001000010000",
									"0001001000010001",
									"0001001000010010",
									"0001001000010011",
									"0001001000010100",
									"0001001000010101",
									"0001001000010110",
									"0001001000010111",
									"0001001000011000",
									"0001001000011001",
									"0001001000100000",
									"0001001000100001",
									"0001001000100010",
									"0001001000100011",
									"0001001000100100",
									"0001001000100101",
									"0001001000100110",
									"0001001000100111",
									"0001001000101000",
									"0001001000101001",
									"0001001000110000",
									"0001001000110001",
									"0001001000110010",
									"0001001000110011",
									"0001001000110100",
									"0001001000110101",
									"0001001000110110",
									"0001001000110111",
									"0001001000111000",
									"0001001000111001",
									"0001001001000000",
									"0001001001000001",
									"0001001001000010",
									"0001001001000011",
									"0001001001000100",
									"0001001001000101",
									"0001001001000110",
									"0001001001000111",
									"0001001001001000",
									"0001001001001001",
									"0001001001010000",
									"0001001001010001",
									"0001001001010010",
									"0001001001010011",
									"0001001001010100",
									"0001001001010101",
									"0001001001010110",
									"0001001001010111",
									"0001001001011000",
									"0001001001011001",
									"0001001001100000",
									"0001001001100001",
									"0001001001100010",
									"0001001001100011",
									"0001001001100100",
									"0001001001100101",
									"0001001001100110",
									"0001001001100111",
									"0001001001101000",
									"0001001001101001",
									"0001001001110000",
									"0001001001110001",
									"0001001001110010",
									"0001001001110011",
									"0001001001110100",
									"0001001001110101",
									"0001001001110110",
									"0001001001110111",
									"0001001001111000",
									"0001001001111001",
									"0001001010000000",
									"0001001010000001",
									"0001001010000010",
									"0001001010000011",
									"0001001010000100",
									"0001001010000101",
									"0001001010000110",
									"0001001010000111",
									"0001001010001000",
									"0001001010001001",
									"0001001010010000",
									"0001001010010001",
									"0001001010010010",
									"0001001010010011",
									"0001001010010100",
									"0001001010010101",
									"0001001010010110",
									"0001001010010111",
									"0001001010011000",
									"0001001010011001",
									"0001001100000000",
									"0001001100000001",
									"0001001100000010",
									"0001001100000011",
									"0001001100000100",
									"0001001100000101",
									"0001001100000110",
									"0001001100000111",
									"0001001100001000",
									"0001001100001001",
									"0001001100010000",
									"0001001100010001",
									"0001001100010010",
									"0001001100010011",
									"0001001100010100",
									"0001001100010101",
									"0001001100010110",
									"0001001100010111",
									"0001001100011000",
									"0001001100011001",
									"0001001100100000",
									"0001001100100001",
									"0001001100100010",
									"0001001100100011",
									"0001001100100100",
									"0001001100100101",
									"0001001100100110",
									"0001001100100111",
									"0001001100101000",
									"0001001100101001",
									"0001001100110000",
									"0001001100110001",
									"0001001100110010",
									"0001001100110011",
									"0001001100110100",
									"0001001100110101",
									"0001001100110110",
									"0001001100110111",
									"0001001100111000",
									"0001001100111001",
									"0001001101000000",
									"0001001101000001",
									"0001001101000010",
									"0001001101000011",
									"0001001101000100",
									"0001001101000101",
									"0001001101000110",
									"0001001101000111",
									"0001001101001000",
									"0001001101001001",
									"0001001101010000",
									"0001001101010001",
									"0001001101010010",
									"0001001101010011",
									"0001001101010100",
									"0001001101010101",
									"0001001101010110",
									"0001001101010111",
									"0001001101011000",
									"0001001101011001",
									"0001001101100000",
									"0001001101100001",
									"0001001101100010",
									"0001001101100011",
									"0001001101100100",
									"0001001101100101",
									"0001001101100110",
									"0001001101100111",
									"0001001101101000",
									"0001001101101001",
									"0001001101110000",
									"0001001101110001",
									"0001001101110010",
									"0001001101110011",
									"0001001101110100",
									"0001001101110101",
									"0001001101110110",
									"0001001101110111",
									"0001001101111000",
									"0001001101111001",
									"0001001110000000",
									"0001001110000001",
									"0001001110000010",
									"0001001110000011",
									"0001001110000100",
									"0001001110000101",
									"0001001110000110",
									"0001001110000111",
									"0001001110001000",
									"0001001110001001",
									"0001001110010000",
									"0001001110010001",
									"0001001110010010",
									"0001001110010011",
									"0001001110010100",
									"0001001110010101",
									"0001001110010110",
									"0001001110010111",
									"0001001110011000",
									"0001001110011001",
									"0001010000000000",
									"0001010000000001",
									"0001010000000010",
									"0001010000000011",
									"0001010000000100",
									"0001010000000101",
									"0001010000000110",
									"0001010000000111",
									"0001010000001000",
									"0001010000001001",
									"0001010000010000",
									"0001010000010001",
									"0001010000010010",
									"0001010000010011",
									"0001010000010100",
									"0001010000010101",
									"0001010000010110",
									"0001010000010111",
									"0001010000011000",
									"0001010000011001",
									"0001010000100000",
									"0001010000100001",
									"0001010000100010",
									"0001010000100011",
									"0001010000100100",
									"0001010000100101",
									"0001010000100110",
									"0001010000100111",
									"0001010000101000",
									"0001010000101001",
									"0001010000110000",
									"0001010000110001",
									"0001010000110010",
									"0001010000110011",
									"0001010000110100",
									"0001010000110101",
									"0001010000110110",
									"0001010000110111",
									"0001010000111000",
									"0001010000111001",
									"0001010001000000",
									"0001010001000001",
									"0001010001000010",
									"0001010001000011",
									"0001010001000100",
									"0001010001000101",
									"0001010001000110",
									"0001010001000111",
									"0001010001001000",
									"0001010001001001",
									"0001010001010000",
									"0001010001010001",
									"0001010001010010",
									"0001010001010011",
									"0001010001010100",
									"0001010001010101",
									"0001010001010110",
									"0001010001010111",
									"0001010001011000",
									"0001010001011001",
									"0001010001100000",
									"0001010001100001",
									"0001010001100010",
									"0001010001100011",
									"0001010001100100",
									"0001010001100101",
									"0001010001100110",
									"0001010001100111",
									"0001010001101000",
									"0001010001101001",
									"0001010001110000",
									"0001010001110001",
									"0001010001110010",
									"0001010001110011",
									"0001010001110100",
									"0001010001110101",
									"0001010001110110",
									"0001010001110111",
									"0001010001111000",
									"0001010001111001",
									"0001010010000000",
									"0001010010000001",
									"0001010010000010",
									"0001010010000011",
									"0001010010000100",
									"0001010010000101",
									"0001010010000110",
									"0001010010000111",
									"0001010010001000",
									"0001010010001001",
									"0001010010010000",
									"0001010010010001",
									"0001010010010010",
									"0001010010010011",
									"0001010010010100",
									"0001010010010101",
									"0001010010010110",
									"0001010010010111",
									"0001010010011000",
									"0001010010011001",
									"0001010100000000",
									"0001010100000001",
									"0001010100000010",
									"0001010100000011",
									"0001010100000100",
									"0001010100000101",
									"0001010100000110",
									"0001010100000111",
									"0001010100001000",
									"0001010100001001",
									"0001010100010000",
									"0001010100010001",
									"0001010100010010",
									"0001010100010011",
									"0001010100010100",
									"0001010100010101",
									"0001010100010110",
									"0001010100010111",
									"0001010100011000",
									"0001010100011001",
									"0001010100100000",
									"0001010100100001",
									"0001010100100010",
									"0001010100100011",
									"0001010100100100",
									"0001010100100101",
									"0001010100100110",
									"0001010100100111",
									"0001010100101000",
									"0001010100101001",
									"0001010100110000",
									"0001010100110001",
									"0001010100110010",
									"0001010100110011",
									"0001010100110100",
									"0001010100110101",
									"0001010100110110",
									"0001010100110111",
									"0001010100111000",
									"0001010100111001",
									"0001010101000000",
									"0001010101000001",
									"0001010101000010",
									"0001010101000011",
									"0001010101000100",
									"0001010101000101",
									"0001010101000110",
									"0001010101000111",
									"0001010101001000",
									"0001010101001001",
									"0001010101010000",
									"0001010101010001",
									"0001010101010010",
									"0001010101010011",
									"0001010101010100",
									"0001010101010101",
									"0001010101010110",
									"0001010101010111",
									"0001010101011000",
									"0001010101011001",
									"0001010101100000",
									"0001010101100001",
									"0001010101100010",
									"0001010101100011",
									"0001010101100100",
									"0001010101100101",
									"0001010101100110",
									"0001010101100111",
									"0001010101101000",
									"0001010101101001",
									"0001010101110000",
									"0001010101110001",
									"0001010101110010",
									"0001010101110011",
									"0001010101110100",
									"0001010101110101",
									"0001010101110110",
									"0001010101110111",
									"0001010101111000",
									"0001010101111001",
									"0001010110000000",
									"0001010110000001",
									"0001010110000010",
									"0001010110000011",
									"0001010110000100",
									"0001010110000101",
									"0001010110000110",
									"0001010110000111",
									"0001010110001000",
									"0001010110001001",
									"0001010110010000",
									"0001010110010001",
									"0001010110010010",
									"0001010110010011",
									"0001010110010100",
									"0001010110010101",
									"0001010110010110",
									"0001010110010111",
									"0001010110011000",
									"0001010110011001",
									"0001011000000000",
									"0001011000000001",
									"0001011000000010",
									"0001011000000011",
									"0001011000000100",
									"0001011000000101",
									"0001011000000110",
									"0001011000000111",
									"0001011000001000",
									"0001011000001001",
									"0001011000010000",
									"0001011000010001",
									"0001011000010010",
									"0001011000010011",
									"0001011000010100",
									"0001011000010101",
									"0001011000010110",
									"0001011000010111",
									"0001011000011000",
									"0001011000011001",
									"0001011000100000",
									"0001011000100001",
									"0001011000100010",
									"0001011000100011",
									"0001011000100100",
									"0001011000100101",
									"0001011000100110",
									"0001011000100111",
									"0001011000101000",
									"0001011000101001",
									"0001011000110000",
									"0001011000110001",
									"0001011000110010",
									"0001011000110011",
									"0001011000110100",
									"0001011000110101",
									"0001011000110110",
									"0001011000110111",
									"0001011000111000",
									"0001011000111001",
									"0001011001000000",
									"0001011001000001",
									"0001011001000010",
									"0001011001000011",
									"0001011001000100",
									"0001011001000101",
									"0001011001000110",
									"0001011001000111",
									"0001011001001000",
									"0001011001001001",
									"0001011001010000",
									"0001011001010001",
									"0001011001010010",
									"0001011001010011",
									"0001011001010100",
									"0001011001010101",
									"0001011001010110",
									"0001011001010111",
									"0001011001011000",
									"0001011001011001",
									"0001011001100000",
									"0001011001100001",
									"0001011001100010",
									"0001011001100011",
									"0001011001100100",
									"0001011001100101",
									"0001011001100110",
									"0001011001100111",
									"0001011001101000",
									"0001011001101001",
									"0001011001110000",
									"0001011001110001",
									"0001011001110010",
									"0001011001110011",
									"0001011001110100",
									"0001011001110101",
									"0001011001110110",
									"0001011001110111",
									"0001011001111000",
									"0001011001111001",
									"0001011010000000",
									"0001011010000001",
									"0001011010000010",
									"0001011010000011",
									"0001011010000100",
									"0001011010000101",
									"0001011010000110",
									"0001011010000111",
									"0001011010001000",
									"0001011010001001",
									"0001011010010000",
									"0001011010010001",
									"0001011010010010",
									"0001011010010011",
									"0001011010010100",
									"0001011010010101",
									"0001011010010110",
									"0001011010010111",
									"0001011010011000",
									"0001011010011001",
									"0001011100000000",
									"0001011100000001",
									"0001011100000010",
									"0001011100000011",
									"0001011100000100",
									"0001011100000101",
									"0001011100000110",
									"0001011100000111",
									"0001011100001000",
									"0001011100001001",
									"0001011100010000",
									"0001011100010001",
									"0001011100010010",
									"0001011100010011",
									"0001011100010100",
									"0001011100010101",
									"0001011100010110",
									"0001011100010111",
									"0001011100011000",
									"0001011100011001",
									"0001011100100000",
									"0001011100100001",
									"0001011100100010",
									"0001011100100011",
									"0001011100100100",
									"0001011100100101",
									"0001011100100110",
									"0001011100100111",
									"0001011100101000",
									"0001011100101001",
									"0001011100110000",
									"0001011100110001",
									"0001011100110010",
									"0001011100110011",
									"0001011100110100",
									"0001011100110101",
									"0001011100110110",
									"0001011100110111",
									"0001011100111000",
									"0001011100111001",
									"0001011101000000",
									"0001011101000001",
									"0001011101000010",
									"0001011101000011",
									"0001011101000100",
									"0001011101000101",
									"0001011101000110",
									"0001011101000111",
									"0001011101001000",
									"0001011101001001",
									"0001011101010000",
									"0001011101010001",
									"0001011101010010",
									"0001011101010011",
									"0001011101010100",
									"0001011101010101",
									"0001011101010110",
									"0001011101010111",
									"0001011101011000",
									"0001011101011001",
									"0001011101100000",
									"0001011101100001",
									"0001011101100010",
									"0001011101100011",
									"0001011101100100",
									"0001011101100101",
									"0001011101100110",
									"0001011101100111",
									"0001011101101000",
									"0001011101101001",
									"0001011101110000",
									"0001011101110001",
									"0001011101110010",
									"0001011101110011",
									"0001011101110100",
									"0001011101110101",
									"0001011101110110",
									"0001011101110111",
									"0001011101111000",
									"0001011101111001",
									"0001011110000000",
									"0001011110000001",
									"0001011110000010",
									"0001011110000011",
									"0001011110000100",
									"0001011110000101",
									"0001011110000110",
									"0001011110000111",
									"0001011110001000",
									"0001011110001001",
									"0001011110010000",
									"0001011110010001",
									"0001011110010010",
									"0001011110010011",
									"0001011110010100",
									"0001011110010101",
									"0001011110010110",
									"0001011110010111",
									"0001011110011000",
									"0001011110011001",
									"0001100000000000",
									"0001100000000001",
									"0001100000000010",
									"0001100000000011",
									"0001100000000100",
									"0001100000000101",
									"0001100000000110",
									"0001100000000111",
									"0001100000001000",
									"0001100000001001",
									"0001100000010000",
									"0001100000010001",
									"0001100000010010",
									"0001100000010011",
									"0001100000010100",
									"0001100000010101",
									"0001100000010110",
									"0001100000010111",
									"0001100000011000",
									"0001100000011001",
									"0001100000100000",
									"0001100000100001",
									"0001100000100010",
									"0001100000100011",
									"0001100000100100",
									"0001100000100101",
									"0001100000100110",
									"0001100000100111",
									"0001100000101000",
									"0001100000101001",
									"0001100000110000",
									"0001100000110001",
									"0001100000110010",
									"0001100000110011",
									"0001100000110100",
									"0001100000110101",
									"0001100000110110",
									"0001100000110111",
									"0001100000111000",
									"0001100000111001",
									"0001100001000000",
									"0001100001000001",
									"0001100001000010",
									"0001100001000011",
									"0001100001000100",
									"0001100001000101",
									"0001100001000110",
									"0001100001000111",
									"0001100001001000",
									"0001100001001001",
									"0001100001010000",
									"0001100001010001",
									"0001100001010010",
									"0001100001010011",
									"0001100001010100",
									"0001100001010101",
									"0001100001010110",
									"0001100001010111",
									"0001100001011000",
									"0001100001011001",
									"0001100001100000",
									"0001100001100001",
									"0001100001100010",
									"0001100001100011",
									"0001100001100100",
									"0001100001100101",
									"0001100001100110",
									"0001100001100111",
									"0001100001101000",
									"0001100001101001",
									"0001100001110000",
									"0001100001110001",
									"0001100001110010",
									"0001100001110011",
									"0001100001110100",
									"0001100001110101",
									"0001100001110110",
									"0001100001110111",
									"0001100001111000",
									"0001100001111001",
									"0001100010000000",
									"0001100010000001",
									"0001100010000010",
									"0001100010000011",
									"0001100010000100",
									"0001100010000101",
									"0001100010000110",
									"0001100010000111",
									"0001100010001000",
									"0001100010001001",
									"0001100010010000",
									"0001100010010001",
									"0001100010010010",
									"0001100010010011",
									"0001100010010100",
									"0001100010010101",
									"0001100010010110",
									"0001100010010111",
									"0001100010011000",
									"0001100010011001",
									"0001100100000000",
									"0001100100000001",
									"0001100100000010",
									"0001100100000011",
									"0001100100000100",
									"0001100100000101",
									"0001100100000110",
									"0001100100000111",
									"0001100100001000",
									"0001100100001001",
									"0001100100010000",
									"0001100100010001",
									"0001100100010010",
									"0001100100010011",
									"0001100100010100",
									"0001100100010101",
									"0001100100010110",
									"0001100100010111",
									"0001100100011000",
									"0001100100011001",
									"0001100100100000",
									"0001100100100001",
									"0001100100100010",
									"0001100100100011",
									"0001100100100100",
									"0001100100100101",
									"0001100100100110",
									"0001100100100111",
									"0001100100101000",
									"0001100100101001",
									"0001100100110000",
									"0001100100110001",
									"0001100100110010",
									"0001100100110011",
									"0001100100110100",
									"0001100100110101",
									"0001100100110110",
									"0001100100110111",
									"0001100100111000",
									"0001100100111001",
									"0001100101000000",
									"0001100101000001",
									"0001100101000010",
									"0001100101000011",
									"0001100101000100",
									"0001100101000101",
									"0001100101000110",
									"0001100101000111",
									"0001100101001000",
									"0001100101001001",
									"0001100101010000",
									"0001100101010001",
									"0001100101010010",
									"0001100101010011",
									"0001100101010100",
									"0001100101010101",
									"0001100101010110",
									"0001100101010111",
									"0001100101011000",
									"0001100101011001",
									"0001100101100000",
									"0001100101100001",
									"0001100101100010",
									"0001100101100011",
									"0001100101100100",
									"0001100101100101",
									"0001100101100110",
									"0001100101100111",
									"0001100101101000",
									"0001100101101001",
									"0001100101110000",
									"0001100101110001",
									"0001100101110010",
									"0001100101110011",
									"0001100101110100",
									"0001100101110101",
									"0001100101110110",
									"0001100101110111",
									"0001100101111000",
									"0001100101111001",
									"0001100110000000",
									"0001100110000001",
									"0001100110000010",
									"0001100110000011",
									"0001100110000100",
									"0001100110000101",
									"0001100110000110",
									"0001100110000111",
									"0001100110001000",
									"0001100110001001",
									"0001100110010000",
									"0001100110010001",
									"0001100110010010",
									"0001100110010011",
									"0001100110010100",
									"0001100110010101",
									"0001100110010110",
									"0001100110010111",
									"0001100110011000",
									"0001100110011001",
									"0010000000000000",
									"0010000000000001",
									"0010000000000010",
									"0010000000000011",
									"0010000000000100",
									"0010000000000101",
									"0010000000000110",
									"0010000000000111",
									"0010000000001000",
									"0010000000001001",
									"0010000000010000",
									"0010000000010001",
									"0010000000010010",
									"0010000000010011",
									"0010000000010100",
									"0010000000010101",
									"0010000000010110",
									"0010000000010111",
									"0010000000011000",
									"0010000000011001",
									"0010000000100000",
									"0010000000100001",
									"0010000000100010",
									"0010000000100011",
									"0010000000100100",
									"0010000000100101",
									"0010000000100110",
									"0010000000100111",
									"0010000000101000",
									"0010000000101001",
									"0010000000110000",
									"0010000000110001",
									"0010000000110010",
									"0010000000110011",
									"0010000000110100",
									"0010000000110101",
									"0010000000110110",
									"0010000000110111",
									"0010000000111000",
									"0010000000111001",
									"0010000001000000",
									"0010000001000001",
									"0010000001000010",
									"0010000001000011",
									"0010000001000100",
									"0010000001000101",
									"0010000001000110",
									"0010000001000111",
									"0010000001001000",
									"0010000001001001",
									"0010000001010000",
									"0010000001010001",
									"0010000001010010",
									"0010000001010011",
									"0010000001010100",
									"0010000001010101",
									"0010000001010110",
									"0010000001010111",
									"0010000001011000",
									"0010000001011001",
									"0010000001100000",
									"0010000001100001",
									"0010000001100010",
									"0010000001100011",
									"0010000001100100",
									"0010000001100101",
									"0010000001100110",
									"0010000001100111",
									"0010000001101000",
									"0010000001101001",
									"0010000001110000",
									"0010000001110001",
									"0010000001110010",
									"0010000001110011",
									"0010000001110100",
									"0010000001110101",
									"0010000001110110",
									"0010000001110111",
									"0010000001111000",
									"0010000001111001",
									"0010000010000000",
									"0010000010000001",
									"0010000010000010",
									"0010000010000011",
									"0010000010000100",
									"0010000010000101",
									"0010000010000110",
									"0010000010000111",
									"0010000010001000",
									"0010000010001001",
									"0010000010010000",
									"0010000010010001",
									"0010000010010010",
									"0010000010010011",
									"0010000010010100",
									"0010000010010101",
									"0010000010010110",
									"0010000010010111",
									"0010000010011000",
									"0010000010011001",
									"0010000100000000",
									"0010000100000001",
									"0010000100000010",
									"0010000100000011",
									"0010000100000100",
									"0010000100000101",
									"0010000100000110",
									"0010000100000111",
									"0010000100001000",
									"0010000100001001",
									"0010000100010000",
									"0010000100010001",
									"0010000100010010",
									"0010000100010011",
									"0010000100010100",
									"0010000100010101",
									"0010000100010110",
									"0010000100010111",
									"0010000100011000",
									"0010000100011001",
									"0010000100100000",
									"0010000100100001",
									"0010000100100010",
									"0010000100100011",
									"0010000100100100",
									"0010000100100101",
									"0010000100100110",
									"0010000100100111",
									"0010000100101000",
									"0010000100101001",
									"0010000100110000",
									"0010000100110001",
									"0010000100110010",
									"0010000100110011",
									"0010000100110100",
									"0010000100110101",
									"0010000100110110",
									"0010000100110111",
									"0010000100111000",
									"0010000100111001",
									"0010000101000000",
									"0010000101000001",
									"0010000101000010",
									"0010000101000011",
									"0010000101000100",
									"0010000101000101",
									"0010000101000110",
									"0010000101000111",
									"0010000101001000",
									"0010000101001001",
									"0010000101010000",
									"0010000101010001",
									"0010000101010010",
									"0010000101010011",
									"0010000101010100",
									"0010000101010101",
									"0010000101010110",
									"0010000101010111",
									"0010000101011000",
									"0010000101011001",
									"0010000101100000",
									"0010000101100001",
									"0010000101100010",
									"0010000101100011",
									"0010000101100100",
									"0010000101100101",
									"0010000101100110",
									"0010000101100111",
									"0010000101101000",
									"0010000101101001",
									"0010000101110000",
									"0010000101110001",
									"0010000101110010",
									"0010000101110011",
									"0010000101110100",
									"0010000101110101",
									"0010000101110110",
									"0010000101110111",
									"0010000101111000",
									"0010000101111001",
									"0010000110000000",
									"0010000110000001",
									"0010000110000010",
									"0010000110000011",
									"0010000110000100",
									"0010000110000101",
									"0010000110000110",
									"0010000110000111",
									"0010000110001000",
									"0010000110001001",
									"0010000110010000",
									"0010000110010001",
									"0010000110010010",
									"0010000110010011",
									"0010000110010100",
									"0010000110010101",
									"0010000110010110",
									"0010000110010111",
									"0010000110011000",
									"0010000110011001",
									"0010001000000000",
									"0010001000000001",
									"0010001000000010",
									"0010001000000011",
									"0010001000000100",
									"0010001000000101",
									"0010001000000110",
									"0010001000000111",
									"0010001000001000",
									"0010001000001001",
									"0010001000010000",
									"0010001000010001",
									"0010001000010010",
									"0010001000010011",
									"0010001000010100",
									"0010001000010101",
									"0010001000010110",
									"0010001000010111",
									"0010001000011000",
									"0010001000011001",
									"0010001000100000",
									"0010001000100001",
									"0010001000100010",
									"0010001000100011",
									"0010001000100100",
									"0010001000100101",
									"0010001000100110",
									"0010001000100111",
									"0010001000101000",
									"0010001000101001",
									"0010001000110000",
									"0010001000110001",
									"0010001000110010",
									"0010001000110011",
									"0010001000110100",
									"0010001000110101",
									"0010001000110110",
									"0010001000110111",
									"0010001000111000",
									"0010001000111001",
									"0010001001000000",
									"0010001001000001",
									"0010001001000010",
									"0010001001000011",
									"0010001001000100",
									"0010001001000101",
									"0010001001000110",
									"0010001001000111",
									"0010001001001000",
									"0010001001001001",
									"0010001001010000",
									"0010001001010001",
									"0010001001010010",
									"0010001001010011",
									"0010001001010100",
									"0010001001010101",
									"0010001001010110",
									"0010001001010111",
									"0010001001011000",
									"0010001001011001",
									"0010001001100000",
									"0010001001100001",
									"0010001001100010",
									"0010001001100011",
									"0010001001100100",
									"0010001001100101",
									"0010001001100110",
									"0010001001100111",
									"0010001001101000",
									"0010001001101001",
									"0010001001110000",
									"0010001001110001",
									"0010001001110010",
									"0010001001110011",
									"0010001001110100",
									"0010001001110101",
									"0010001001110110",
									"0010001001110111",
									"0010001001111000",
									"0010001001111001",
									"0010001010000000",
									"0010001010000001",
									"0010001010000010",
									"0010001010000011",
									"0010001010000100",
									"0010001010000101",
									"0010001010000110",
									"0010001010000111",
									"0010001010001000",
									"0010001010001001",
									"0010001010010000",
									"0010001010010001",
									"0010001010010010",
									"0010001010010011",
									"0010001010010100",
									"0010001010010101",
									"0010001010010110",
									"0010001010010111",
									"0010001010011000",
									"0010001010011001",
									"0010001100000000",
									"0010001100000001",
									"0010001100000010",
									"0010001100000011",
									"0010001100000100",
									"0010001100000101",
									"0010001100000110",
									"0010001100000111",
									"0010001100001000",
									"0010001100001001",
									"0010001100010000",
									"0010001100010001",
									"0010001100010010",
									"0010001100010011",
									"0010001100010100",
									"0010001100010101",
									"0010001100010110",
									"0010001100010111",
									"0010001100011000",
									"0010001100011001",
									"0010001100100000",
									"0010001100100001",
									"0010001100100010",
									"0010001100100011",
									"0010001100100100",
									"0010001100100101",
									"0010001100100110",
									"0010001100100111",
									"0010001100101000",
									"0010001100101001",
									"0010001100110000",
									"0010001100110001",
									"0010001100110010",
									"0010001100110011",
									"0010001100110100",
									"0010001100110101",
									"0010001100110110",
									"0010001100110111",
									"0010001100111000",
									"0010001100111001",
									"0010001101000000",
									"0010001101000001",
									"0010001101000010",
									"0010001101000011",
									"0010001101000100",
									"0010001101000101",
									"0010001101000110",
									"0010001101000111",
									"0010001101001000",
									"0010001101001001",
									"0010001101010000",
									"0010001101010001",
									"0010001101010010",
									"0010001101010011",
									"0010001101010100",
									"0010001101010101",
									"0010001101010110",
									"0010001101010111",
									"0010001101011000",
									"0010001101011001",
									"0010001101100000",
									"0010001101100001",
									"0010001101100010",
									"0010001101100011",
									"0010001101100100",
									"0010001101100101",
									"0010001101100110",
									"0010001101100111",
									"0010001101101000",
									"0010001101101001",
									"0010001101110000",
									"0010001101110001",
									"0010001101110010",
									"0010001101110011",
									"0010001101110100",
									"0010001101110101",
									"0010001101110110",
									"0010001101110111",
									"0010001101111000",
									"0010001101111001",
									"0010001110000000",
									"0010001110000001",
									"0010001110000010",
									"0010001110000011",
									"0010001110000100",
									"0010001110000101",
									"0010001110000110",
									"0010001110000111",
									"0010001110001000",
									"0010001110001001",
									"0010001110010000",
									"0010001110010001",
									"0010001110010010",
									"0010001110010011",
									"0010001110010100",
									"0010001110010101",
									"0010001110010110",
									"0010001110010111",
									"0010001110011000",
									"0010001110011001",
									"0010010000000000",
									"0010010000000001",
									"0010010000000010",
									"0010010000000011",
									"0010010000000100",
									"0010010000000101",
									"0010010000000110",
									"0010010000000111",
									"0010010000001000",
									"0010010000001001",
									"0010010000010000",
									"0010010000010001",
									"0010010000010010",
									"0010010000010011",
									"0010010000010100",
									"0010010000010101",
									"0010010000010110",
									"0010010000010111",
									"0010010000011000",
									"0010010000011001",
									"0010010000100000",
									"0010010000100001",
									"0010010000100010",
									"0010010000100011",
									"0010010000100100",
									"0010010000100101",
									"0010010000100110",
									"0010010000100111",
									"0010010000101000",
									"0010010000101001",
									"0010010000110000",
									"0010010000110001",
									"0010010000110010",
									"0010010000110011",
									"0010010000110100",
									"0010010000110101",
									"0010010000110110",
									"0010010000110111",
									"0010010000111000",
									"0010010000111001",
									"0010010001000000",
									"0010010001000001",
									"0010010001000010",
									"0010010001000011",
									"0010010001000100",
									"0010010001000101",
									"0010010001000110",
									"0010010001000111",
									"0010010001001000",
									"0010010001001001",
									"0010010001010000",
									"0010010001010001",
									"0010010001010010",
									"0010010001010011",
									"0010010001010100",
									"0010010001010101",
									"0010010001010110",
									"0010010001010111",
									"0010010001011000",
									"0010010001011001",
									"0010010001100000",
									"0010010001100001",
									"0010010001100010",
									"0010010001100011",
									"0010010001100100",
									"0010010001100101",
									"0010010001100110",
									"0010010001100111",
									"0010010001101000",
									"0010010001101001",
									"0010010001110000",
									"0010010001110001",
									"0010010001110010",
									"0010010001110011",
									"0010010001110100",
									"0010010001110101",
									"0010010001110110",
									"0010010001110111",
									"0010010001111000",
									"0010010001111001",
									"0010010010000000",
									"0010010010000001",
									"0010010010000010",
									"0010010010000011",
									"0010010010000100",
									"0010010010000101",
									"0010010010000110",
									"0010010010000111",
									"0010010010001000",
									"0010010010001001",
									"0010010010010000",
									"0010010010010001",
									"0010010010010010",
									"0010010010010011",
									"0010010010010100",
									"0010010010010101",
									"0010010010010110",
									"0010010010010111",
									"0010010010011000",
									"0010010010011001",
									"0010010100000000",
									"0010010100000001",
									"0010010100000010",
									"0010010100000011",
									"0010010100000100",
									"0010010100000101",
									"0010010100000110",
									"0010010100000111",
									"0010010100001000",
									"0010010100001001",
									"0010010100010000",
									"0010010100010001",
									"0010010100010010",
									"0010010100010011",
									"0010010100010100",
									"0010010100010101",
									"0010010100010110",
									"0010010100010111",
									"0010010100011000",
									"0010010100011001",
									"0010010100100000",
									"0010010100100001",
									"0010010100100010",
									"0010010100100011",
									"0010010100100100",
									"0010010100100101",
									"0010010100100110",
									"0010010100100111",
									"0010010100101000",
									"0010010100101001",
									"0010010100110000",
									"0010010100110001",
									"0010010100110010",
									"0010010100110011",
									"0010010100110100",
									"0010010100110101",
									"0010010100110110",
									"0010010100110111",
									"0010010100111000",
									"0010010100111001",
									"0010010101000000",
									"0010010101000001",
									"0010010101000010",
									"0010010101000011",
									"0010010101000100",
									"0010010101000101",
									"0010010101000110",
									"0010010101000111",
									"0010010101001000",
									"0010010101001001",
									"0010010101010000",
									"0010010101010001",
									"0010010101010010",
									"0010010101010011",
									"0010010101010100",
									"0010010101010101",
									"0010010101010110",
									"0010010101010111",
									"0010010101011000",
									"0010010101011001",
									"0010010101100000",
									"0010010101100001",
									"0010010101100010",
									"0010010101100011",
									"0010010101100100",
									"0010010101100101",
									"0010010101100110",
									"0010010101100111",
									"0010010101101000",
									"0010010101101001",
									"0010010101110000",
									"0010010101110001",
									"0010010101110010",
									"0010010101110011",
									"0010010101110100",
									"0010010101110101",
									"0010010101110110",
									"0010010101110111",
									"0010010101111000",
									"0010010101111001",
									"0010010110000000",
									"0010010110000001",
									"0010010110000010",
									"0010010110000011",
									"0010010110000100",
									"0010010110000101",
									"0010010110000110",
									"0010010110000111",
									"0010010110001000",
									"0010010110001001",
									"0010010110010000",
									"0010010110010001",
									"0010010110010010",
									"0010010110010011",
									"0010010110010100",
									"0010010110010101",
									"0010010110010110",
									"0010010110010111",
									"0010010110011000",
									"0010010110011001",
									"0010011000000000",
									"0010011000000001",
									"0010011000000010",
									"0010011000000011",
									"0010011000000100",
									"0010011000000101",
									"0010011000000110",
									"0010011000000111",
									"0010011000001000",
									"0010011000001001",
									"0010011000010000",
									"0010011000010001",
									"0010011000010010",
									"0010011000010011",
									"0010011000010100",
									"0010011000010101",
									"0010011000010110",
									"0010011000010111",
									"0010011000011000",
									"0010011000011001",
									"0010011000100000",
									"0010011000100001",
									"0010011000100010",
									"0010011000100011",
									"0010011000100100",
									"0010011000100101",
									"0010011000100110",
									"0010011000100111",
									"0010011000101000",
									"0010011000101001",
									"0010011000110000",
									"0010011000110001",
									"0010011000110010",
									"0010011000110011",
									"0010011000110100",
									"0010011000110101",
									"0010011000110110",
									"0010011000110111",
									"0010011000111000",
									"0010011000111001",
									"0010011001000000",
									"0010011001000001",
									"0010011001000010",
									"0010011001000011",
									"0010011001000100",
									"0010011001000101",
									"0010011001000110",
									"0010011001000111",
									"0010011001001000",
									"0010011001001001",
									"0010011001010000",
									"0010011001010001",
									"0010011001010010",
									"0010011001010011",
									"0010011001010100",
									"0010011001010101",
									"0010011001010110",
									"0010011001010111",
									"0010011001011000",
									"0010011001011001",
									"0010011001100000",
									"0010011001100001",
									"0010011001100010",
									"0010011001100011",
									"0010011001100100",
									"0010011001100101",
									"0010011001100110",
									"0010011001100111",
									"0010011001101000",
									"0010011001101001",
									"0010011001110000",
									"0010011001110001",
									"0010011001110010",
									"0010011001110011",
									"0010011001110100",
									"0010011001110101",
									"0010011001110110",
									"0010011001110111",
									"0010011001111000",
									"0010011001111001",
									"0010011010000000",
									"0010011010000001",
									"0010011010000010",
									"0010011010000011",
									"0010011010000100",
									"0010011010000101",
									"0010011010000110",
									"0010011010000111",
									"0010011010001000",
									"0010011010001001",
									"0010011010010000",
									"0010011010010001",
									"0010011010010010",
									"0010011010010011",
									"0010011010010100",
									"0010011010010101",
									"0010011010010110",
									"0010011010010111",
									"0010011010011000",
									"0010011010011001",
									"0010011100000000",
									"0010011100000001",
									"0010011100000010",
									"0010011100000011",
									"0010011100000100",
									"0010011100000101",
									"0010011100000110",
									"0010011100000111",
									"0010011100001000",
									"0010011100001001",
									"0010011100010000",
									"0010011100010001",
									"0010011100010010",
									"0010011100010011",
									"0010011100010100",
									"0010011100010101",
									"0010011100010110",
									"0010011100010111",
									"0010011100011000",
									"0010011100011001",
									"0010011100100000",
									"0010011100100001",
									"0010011100100010",
									"0010011100100011",
									"0010011100100100",
									"0010011100100101",
									"0010011100100110",
									"0010011100100111",
									"0010011100101000",
									"0010011100101001",
									"0010011100110000",
									"0010011100110001",
									"0010011100110010",
									"0010011100110011",
									"0010011100110100",
									"0010011100110101",
									"0010011100110110",
									"0010011100110111",
									"0010011100111000",
									"0010011100111001",
									"0010011101000000",
									"0010011101000001",
									"0010011101000010",
									"0010011101000011",
									"0010011101000100",
									"0010011101000101",
									"0010011101000110",
									"0010011101000111",
									"0010011101001000",
									"0010011101001001",
									"0010011101010000",
									"0010011101010001",
									"0010011101010010",
									"0010011101010011",
									"0010011101010100",
									"0010011101010101",
									"0010011101010110",
									"0010011101010111",
									"0010011101011000",
									"0010011101011001",
									"0010011101100000",
									"0010011101100001",
									"0010011101100010",
									"0010011101100011",
									"0010011101100100",
									"0010011101100101",
									"0010011101100110",
									"0010011101100111",
									"0010011101101000",
									"0010011101101001",
									"0010011101110000",
									"0010011101110001",
									"0010011101110010",
									"0010011101110011",
									"0010011101110100",
									"0010011101110101",
									"0010011101110110",
									"0010011101110111",
									"0010011101111000",
									"0010011101111001",
									"0010011110000000",
									"0010011110000001",
									"0010011110000010",
									"0010011110000011",
									"0010011110000100",
									"0010011110000101",
									"0010011110000110",
									"0010011110000111",
									"0010011110001000",
									"0010011110001001",
									"0010011110010000",
									"0010011110010001",
									"0010011110010010",
									"0010011110010011",
									"0010011110010100",
									"0010011110010101",
									"0010011110010110",
									"0010011110010111",
									"0010011110011000",
									"0010011110011001",
									"0010100000000000",
									"0010100000000001",
									"0010100000000010",
									"0010100000000011",
									"0010100000000100",
									"0010100000000101",
									"0010100000000110",
									"0010100000000111",
									"0010100000001000",
									"0010100000001001",
									"0010100000010000",
									"0010100000010001",
									"0010100000010010",
									"0010100000010011",
									"0010100000010100",
									"0010100000010101",
									"0010100000010110",
									"0010100000010111",
									"0010100000011000",
									"0010100000011001",
									"0010100000100000",
									"0010100000100001",
									"0010100000100010",
									"0010100000100011",
									"0010100000100100",
									"0010100000100101",
									"0010100000100110",
									"0010100000100111",
									"0010100000101000",
									"0010100000101001",
									"0010100000110000",
									"0010100000110001",
									"0010100000110010",
									"0010100000110011",
									"0010100000110100",
									"0010100000110101",
									"0010100000110110",
									"0010100000110111",
									"0010100000111000",
									"0010100000111001",
									"0010100001000000",
									"0010100001000001",
									"0010100001000010",
									"0010100001000011",
									"0010100001000100",
									"0010100001000101",
									"0010100001000110",
									"0010100001000111",
									"0010100001001000",
									"0010100001001001",
									"0010100001010000",
									"0010100001010001",
									"0010100001010010",
									"0010100001010011",
									"0010100001010100",
									"0010100001010101",
									"0010100001010110",
									"0010100001010111",
									"0010100001011000",
									"0010100001011001",
									"0010100001100000",
									"0010100001100001",
									"0010100001100010",
									"0010100001100011",
									"0010100001100100",
									"0010100001100101",
									"0010100001100110",
									"0010100001100111",
									"0010100001101000",
									"0010100001101001",
									"0010100001110000",
									"0010100001110001",
									"0010100001110010",
									"0010100001110011",
									"0010100001110100",
									"0010100001110101",
									"0010100001110110",
									"0010100001110111",
									"0010100001111000",
									"0010100001111001",
									"0010100010000000",
									"0010100010000001",
									"0010100010000010",
									"0010100010000011",
									"0010100010000100",
									"0010100010000101",
									"0010100010000110",
									"0010100010000111",
									"0010100010001000",
									"0010100010001001",
									"0010100010010000",
									"0010100010010001",
									"0010100010010010",
									"0010100010010011",
									"0010100010010100",
									"0010100010010101",
									"0010100010010110",
									"0010100010010111",
									"0010100010011000",
									"0010100010011001",
									"0010100100000000",
									"0010100100000001",
									"0010100100000010",
									"0010100100000011",
									"0010100100000100",
									"0010100100000101",
									"0010100100000110",
									"0010100100000111",
									"0010100100001000",
									"0010100100001001",
									"0010100100010000",
									"0010100100010001",
									"0010100100010010",
									"0010100100010011",
									"0010100100010100",
									"0010100100010101",
									"0010100100010110",
									"0010100100010111",
									"0010100100011000",
									"0010100100011001",
									"0010100100100000",
									"0010100100100001",
									"0010100100100010",
									"0010100100100011",
									"0010100100100100",
									"0010100100100101",
									"0010100100100110",
									"0010100100100111",
									"0010100100101000",
									"0010100100101001",
									"0010100100110000",
									"0010100100110001",
									"0010100100110010",
									"0010100100110011",
									"0010100100110100",
									"0010100100110101",
									"0010100100110110",
									"0010100100110111",
									"0010100100111000",
									"0010100100111001",
									"0010100101000000",
									"0010100101000001",
									"0010100101000010",
									"0010100101000011",
									"0010100101000100",
									"0010100101000101",
									"0010100101000110",
									"0010100101000111",
									"0010100101001000",
									"0010100101001001",
									"0010100101010000",
									"0010100101010001",
									"0010100101010010",
									"0010100101010011",
									"0010100101010100",
									"0010100101010101",
									"0010100101010110",
									"0010100101010111",
									"0010100101011000",
									"0010100101011001",
									"0010100101100000",
									"0010100101100001",
									"0010100101100010",
									"0010100101100011",
									"0010100101100100",
									"0010100101100101",
									"0010100101100110",
									"0010100101100111",
									"0010100101101000",
									"0010100101101001",
									"0010100101110000",
									"0010100101110001",
									"0010100101110010",
									"0010100101110011",
									"0010100101110100",
									"0010100101110101",
									"0010100101110110",
									"0010100101110111",
									"0010100101111000",
									"0010100101111001",
									"0010100110000000",
									"0010100110000001",
									"0010100110000010",
									"0010100110000011",
									"0010100110000100",
									"0010100110000101",
									"0010100110000110",
									"0010100110000111",
									"0010100110001000",
									"0010100110001001",
									"0010100110010000",
									"0010100110010001",
									"0010100110010010",
									"0010100110010011",
									"0010100110010100",
									"0010100110010101",
									"0010100110010110",
									"0010100110010111",
									"0010100110011000",
									"0010100110011001",
									"0011000000000000",
									"0011000000000001",
									"0011000000000010",
									"0011000000000011",
									"0011000000000100",
									"0011000000000101",
									"0011000000000110",
									"0011000000000111",
									"0011000000001000",
									"0011000000001001",
									"0011000000010000",
									"0011000000010001",
									"0011000000010010",
									"0011000000010011",
									"0011000000010100",
									"0011000000010101",
									"0011000000010110",
									"0011000000010111",
									"0011000000011000",
									"0011000000011001",
									"0011000000100000",
									"0011000000100001",
									"0011000000100010",
									"0011000000100011",
									"0011000000100100",
									"0011000000100101",
									"0011000000100110",
									"0011000000100111",
									"0011000000101000",
									"0011000000101001",
									"0011000000110000",
									"0011000000110001",
									"0011000000110010",
									"0011000000110011",
									"0011000000110100",
									"0011000000110101",
									"0011000000110110",
									"0011000000110111",
									"0011000000111000",
									"0011000000111001",
									"0011000001000000",
									"0011000001000001",
									"0011000001000010",
									"0011000001000011",
									"0011000001000100",
									"0011000001000101",
									"0011000001000110",
									"0011000001000111",
									"0011000001001000",
									"0011000001001001",
									"0011000001010000",
									"0011000001010001",
									"0011000001010010",
									"0011000001010011",
									"0011000001010100",
									"0011000001010101",
									"0011000001010110",
									"0011000001010111",
									"0011000001011000",
									"0011000001011001",
									"0011000001100000",
									"0011000001100001",
									"0011000001100010",
									"0011000001100011",
									"0011000001100100",
									"0011000001100101",
									"0011000001100110",
									"0011000001100111",
									"0011000001101000",
									"0011000001101001",
									"0011000001110000",
									"0011000001110001",
									"0011000001110010",
									"0011000001110011",
									"0011000001110100",
									"0011000001110101",
									"0011000001110110",
									"0011000001110111",
									"0011000001111000",
									"0011000001111001",
									"0011000010000000",
									"0011000010000001",
									"0011000010000010",
									"0011000010000011",
									"0011000010000100",
									"0011000010000101",
									"0011000010000110",
									"0011000010000111",
									"0011000010001000",
									"0011000010001001",
									"0011000010010000",
									"0011000010010001",
									"0011000010010010",
									"0011000010010011",
									"0011000010010100",
									"0011000010010101",
									"0011000010010110",
									"0011000010010111",
									"0011000010011000",
									"0011000010011001",
									"0011000100000000",
									"0011000100000001",
									"0011000100000010",
									"0011000100000011",
									"0011000100000100",
									"0011000100000101",
									"0011000100000110",
									"0011000100000111",
									"0011000100001000",
									"0011000100001001",
									"0011000100010000",
									"0011000100010001",
									"0011000100010010",
									"0011000100010011",
									"0011000100010100",
									"0011000100010101",
									"0011000100010110",
									"0011000100010111",
									"0011000100011000",
									"0011000100011001",
									"0011000100100000",
									"0011000100100001",
									"0011000100100010",
									"0011000100100011",
									"0011000100100100",
									"0011000100100101",
									"0011000100100110",
									"0011000100100111",
									"0011000100101000",
									"0011000100101001",
									"0011000100110000",
									"0011000100110001",
									"0011000100110010",
									"0011000100110011",
									"0011000100110100",
									"0011000100110101",
									"0011000100110110",
									"0011000100110111",
									"0011000100111000",
									"0011000100111001",
									"0011000101000000",
									"0011000101000001",
									"0011000101000010",
									"0011000101000011",
									"0011000101000100",
									"0011000101000101",
									"0011000101000110",
									"0011000101000111",
									"0011000101001000",
									"0011000101001001",
									"0011000101010000",
									"0011000101010001",
									"0011000101010010",
									"0011000101010011",
									"0011000101010100",
									"0011000101010101",
									"0011000101010110",
									"0011000101010111",
									"0011000101011000",
									"0011000101011001",
									"0011000101100000",
									"0011000101100001",
									"0011000101100010",
									"0011000101100011",
									"0011000101100100",
									"0011000101100101",
									"0011000101100110",
									"0011000101100111",
									"0011000101101000",
									"0011000101101001",
									"0011000101110000",
									"0011000101110001",
									"0011000101110010",
									"0011000101110011",
									"0011000101110100",
									"0011000101110101",
									"0011000101110110",
									"0011000101110111",
									"0011000101111000",
									"0011000101111001",
									"0011000110000000",
									"0011000110000001",
									"0011000110000010",
									"0011000110000011",
									"0011000110000100",
									"0011000110000101",
									"0011000110000110",
									"0011000110000111",
									"0011000110001000",
									"0011000110001001",
									"0011000110010000",
									"0011000110010001",
									"0011000110010010",
									"0011000110010011",
									"0011000110010100",
									"0011000110010101",
									"0011000110010110",
									"0011000110010111",
									"0011000110011000",
									"0011000110011001",
									"0011001000000000",
									"0011001000000001",
									"0011001000000010",
									"0011001000000011",
									"0011001000000100",
									"0011001000000101",
									"0011001000000110",
									"0011001000000111",
									"0011001000001000",
									"0011001000001001",
									"0011001000010000",
									"0011001000010001",
									"0011001000010010",
									"0011001000010011",
									"0011001000010100",
									"0011001000010101",
									"0011001000010110",
									"0011001000010111",
									"0011001000011000",
									"0011001000011001",
									"0011001000100000",
									"0011001000100001",
									"0011001000100010",
									"0011001000100011",
									"0011001000100100",
									"0011001000100101",
									"0011001000100110",
									"0011001000100111",
									"0011001000101000",
									"0011001000101001",
									"0011001000110000",
									"0011001000110001",
									"0011001000110010",
									"0011001000110011",
									"0011001000110100",
									"0011001000110101",
									"0011001000110110",
									"0011001000110111",
									"0011001000111000",
									"0011001000111001",
									"0011001001000000",
									"0011001001000001",
									"0011001001000010",
									"0011001001000011",
									"0011001001000100",
									"0011001001000101",
									"0011001001000110",
									"0011001001000111",
									"0011001001001000",
									"0011001001001001",
									"0011001001010000",
									"0011001001010001",
									"0011001001010010",
									"0011001001010011",
									"0011001001010100",
									"0011001001010101",
									"0011001001010110",
									"0011001001010111",
									"0011001001011000",
									"0011001001011001",
									"0011001001100000",
									"0011001001100001",
									"0011001001100010",
									"0011001001100011",
									"0011001001100100",
									"0011001001100101",
									"0011001001100110",
									"0011001001100111",
									"0011001001101000",
									"0011001001101001",
									"0011001001110000",
									"0011001001110001",
									"0011001001110010",
									"0011001001110011",
									"0011001001110100",
									"0011001001110101",
									"0011001001110110",
									"0011001001110111",
									"0011001001111000",
									"0011001001111001",
									"0011001010000000",
									"0011001010000001",
									"0011001010000010",
									"0011001010000011",
									"0011001010000100",
									"0011001010000101",
									"0011001010000110",
									"0011001010000111",
									"0011001010001000",
									"0011001010001001",
									"0011001010010000",
									"0011001010010001",
									"0011001010010010",
									"0011001010010011",
									"0011001010010100",
									"0011001010010101",
									"0011001010010110",
									"0011001010010111",
									"0011001010011000",
									"0011001010011001",
									"0011001100000000",
									"0011001100000001",
									"0011001100000010",
									"0011001100000011",
									"0011001100000100",
									"0011001100000101",
									"0011001100000110",
									"0011001100000111",
									"0011001100001000",
									"0011001100001001",
									"0011001100010000",
									"0011001100010001",
									"0011001100010010",
									"0011001100010011",
									"0011001100010100",
									"0011001100010101",
									"0011001100010110",
									"0011001100010111",
									"0011001100011000",
									"0011001100011001",
									"0011001100100000",
									"0011001100100001",
									"0011001100100010",
									"0011001100100011",
									"0011001100100100",
									"0011001100100101",
									"0011001100100110",
									"0011001100100111",
									"0011001100101000",
									"0011001100101001",
									"0011001100110000",
									"0011001100110001",
									"0011001100110010",
									"0011001100110011",
									"0011001100110100",
									"0011001100110101",
									"0011001100110110",
									"0011001100110111",
									"0011001100111000",
									"0011001100111001",
									"0011001101000000",
									"0011001101000001",
									"0011001101000010",
									"0011001101000011",
									"0011001101000100",
									"0011001101000101",
									"0011001101000110",
									"0011001101000111",
									"0011001101001000",
									"0011001101001001",
									"0011001101010000",
									"0011001101010001",
									"0011001101010010",
									"0011001101010011",
									"0011001101010100",
									"0011001101010101",
									"0011001101010110",
									"0011001101010111",
									"0011001101011000",
									"0011001101011001",
									"0011001101100000",
									"0011001101100001",
									"0011001101100010",
									"0011001101100011",
									"0011001101100100",
									"0011001101100101",
									"0011001101100110",
									"0011001101100111",
									"0011001101101000",
									"0011001101101001",
									"0011001101110000",
									"0011001101110001",
									"0011001101110010",
									"0011001101110011",
									"0011001101110100",
									"0011001101110101",
									"0011001101110110",
									"0011001101110111",
									"0011001101111000",
									"0011001101111001",
									"0011001110000000",
									"0011001110000001",
									"0011001110000010",
									"0011001110000011",
									"0011001110000100",
									"0011001110000101",
									"0011001110000110",
									"0011001110000111",
									"0011001110001000",
									"0011001110001001",
									"0011001110010000",
									"0011001110010001",
									"0011001110010010",
									"0011001110010011",
									"0011001110010100",
									"0011001110010101",
									"0011001110010110",
									"0011001110010111",
									"0011001110011000",
									"0011001110011001",
									"0011010000000000",
									"0011010000000001",
									"0011010000000010",
									"0011010000000011",
									"0011010000000100",
									"0011010000000101",
									"0011010000000110",
									"0011010000000111",
									"0011010000001000",
									"0011010000001001",
									"0011010000010000",
									"0011010000010001",
									"0011010000010010",
									"0011010000010011",
									"0011010000010100",
									"0011010000010101",
									"0011010000010110",
									"0011010000010111",
									"0011010000011000",
									"0011010000011001",
									"0011010000100000",
									"0011010000100001",
									"0011010000100010",
									"0011010000100011",
									"0011010000100100",
									"0011010000100101",
									"0011010000100110",
									"0011010000100111",
									"0011010000101000",
									"0011010000101001",
									"0011010000110000",
									"0011010000110001",
									"0011010000110010",
									"0011010000110011",
									"0011010000110100",
									"0011010000110101",
									"0011010000110110",
									"0011010000110111",
									"0011010000111000",
									"0011010000111001",
									"0011010001000000",
									"0011010001000001",
									"0011010001000010",
									"0011010001000011",
									"0011010001000100",
									"0011010001000101",
									"0011010001000110",
									"0011010001000111",
									"0011010001001000",
									"0011010001001001",
									"0011010001010000",
									"0011010001010001",
									"0011010001010010",
									"0011010001010011",
									"0011010001010100",
									"0011010001010101",
									"0011010001010110",
									"0011010001010111",
									"0011010001011000",
									"0011010001011001",
									"0011010001100000",
									"0011010001100001",
									"0011010001100010",
									"0011010001100011",
									"0011010001100100",
									"0011010001100101",
									"0011010001100110",
									"0011010001100111",
									"0011010001101000",
									"0011010001101001",
									"0011010001110000",
									"0011010001110001",
									"0011010001110010",
									"0011010001110011",
									"0011010001110100",
									"0011010001110101",
									"0011010001110110",
									"0011010001110111",
									"0011010001111000",
									"0011010001111001",
									"0011010010000000",
									"0011010010000001",
									"0011010010000010",
									"0011010010000011",
									"0011010010000100",
									"0011010010000101",
									"0011010010000110",
									"0011010010000111",
									"0011010010001000",
									"0011010010001001",
									"0011010010010000",
									"0011010010010001",
									"0011010010010010",
									"0011010010010011",
									"0011010010010100",
									"0011010010010101",
									"0011010010010110",
									"0011010010010111",
									"0011010010011000",
									"0011010010011001",
									"0011010100000000",
									"0011010100000001",
									"0011010100000010",
									"0011010100000011",
									"0011010100000100",
									"0011010100000101",
									"0011010100000110",
									"0011010100000111",
									"0011010100001000",
									"0011010100001001",
									"0011010100010000",
									"0011010100010001",
									"0011010100010010",
									"0011010100010011",
									"0011010100010100",
									"0011010100010101",
									"0011010100010110",
									"0011010100010111",
									"0011010100011000",
									"0011010100011001",
									"0011010100100000",
									"0011010100100001",
									"0011010100100010",
									"0011010100100011",
									"0011010100100100",
									"0011010100100101",
									"0011010100100110",
									"0011010100100111",
									"0011010100101000",
									"0011010100101001",
									"0011010100110000",
									"0011010100110001",
									"0011010100110010",
									"0011010100110011",
									"0011010100110100",
									"0011010100110101",
									"0011010100110110",
									"0011010100110111",
									"0011010100111000",
									"0011010100111001",
									"0011010101000000",
									"0011010101000001",
									"0011010101000010",
									"0011010101000011",
									"0011010101000100",
									"0011010101000101",
									"0011010101000110",
									"0011010101000111",
									"0011010101001000",
									"0011010101001001",
									"0011010101010000",
									"0011010101010001",
									"0011010101010010",
									"0011010101010011",
									"0011010101010100",
									"0011010101010101",
									"0011010101010110",
									"0011010101010111",
									"0011010101011000",
									"0011010101011001",
									"0011010101100000",
									"0011010101100001",
									"0011010101100010",
									"0011010101100011",
									"0011010101100100",
									"0011010101100101",
									"0011010101100110",
									"0011010101100111",
									"0011010101101000",
									"0011010101101001",
									"0011010101110000",
									"0011010101110001",
									"0011010101110010",
									"0011010101110011",
									"0011010101110100",
									"0011010101110101",
									"0011010101110110",
									"0011010101110111",
									"0011010101111000",
									"0011010101111001",
									"0011010110000000",
									"0011010110000001",
									"0011010110000010",
									"0011010110000011",
									"0011010110000100",
									"0011010110000101",
									"0011010110000110",
									"0011010110000111",
									"0011010110001000",
									"0011010110001001",
									"0011010110010000",
									"0011010110010001",
									"0011010110010010",
									"0011010110010011",
									"0011010110010100",
									"0011010110010101",
									"0011010110010110",
									"0011010110010111",
									"0011010110011000",
									"0011010110011001",
									"0011011000000000",
									"0011011000000001",
									"0011011000000010",
									"0011011000000011",
									"0011011000000100",
									"0011011000000101",
									"0011011000000110",
									"0011011000000111",
									"0011011000001000",
									"0011011000001001",
									"0011011000010000",
									"0011011000010001",
									"0011011000010010",
									"0011011000010011",
									"0011011000010100",
									"0011011000010101",
									"0011011000010110",
									"0011011000010111",
									"0011011000011000",
									"0011011000011001",
									"0011011000100000",
									"0011011000100001",
									"0011011000100010",
									"0011011000100011",
									"0011011000100100",
									"0011011000100101",
									"0011011000100110",
									"0011011000100111",
									"0011011000101000",
									"0011011000101001",
									"0011011000110000",
									"0011011000110001",
									"0011011000110010",
									"0011011000110011",
									"0011011000110100",
									"0011011000110101",
									"0011011000110110",
									"0011011000110111",
									"0011011000111000",
									"0011011000111001",
									"0011011001000000",
									"0011011001000001",
									"0011011001000010",
									"0011011001000011",
									"0011011001000100",
									"0011011001000101",
									"0011011001000110",
									"0011011001000111",
									"0011011001001000",
									"0011011001001001",
									"0011011001010000",
									"0011011001010001",
									"0011011001010010",
									"0011011001010011",
									"0011011001010100",
									"0011011001010101",
									"0011011001010110",
									"0011011001010111",
									"0011011001011000",
									"0011011001011001",
									"0011011001100000",
									"0011011001100001",
									"0011011001100010",
									"0011011001100011",
									"0011011001100100",
									"0011011001100101",
									"0011011001100110",
									"0011011001100111",
									"0011011001101000",
									"0011011001101001",
									"0011011001110000",
									"0011011001110001",
									"0011011001110010",
									"0011011001110011",
									"0011011001110100",
									"0011011001110101",
									"0011011001110110",
									"0011011001110111",
									"0011011001111000",
									"0011011001111001",
									"0011011010000000",
									"0011011010000001",
									"0011011010000010",
									"0011011010000011",
									"0011011010000100",
									"0011011010000101",
									"0011011010000110",
									"0011011010000111",
									"0011011010001000",
									"0011011010001001",
									"0011011010010000",
									"0011011010010001",
									"0011011010010010",
									"0011011010010011",
									"0011011010010100",
									"0011011010010101",
									"0011011010010110",
									"0011011010010111",
									"0011011010011000",
									"0011011010011001",
									"0011011100000000",
									"0011011100000001",
									"0011011100000010",
									"0011011100000011",
									"0011011100000100",
									"0011011100000101",
									"0011011100000110",
									"0011011100000111",
									"0011011100001000",
									"0011011100001001",
									"0011011100010000",
									"0011011100010001",
									"0011011100010010",
									"0011011100010011",
									"0011011100010100",
									"0011011100010101",
									"0011011100010110",
									"0011011100010111",
									"0011011100011000",
									"0011011100011001",
									"0011011100100000",
									"0011011100100001",
									"0011011100100010",
									"0011011100100011",
									"0011011100100100",
									"0011011100100101",
									"0011011100100110",
									"0011011100100111",
									"0011011100101000",
									"0011011100101001",
									"0011011100110000",
									"0011011100110001",
									"0011011100110010",
									"0011011100110011",
									"0011011100110100",
									"0011011100110101",
									"0011011100110110",
									"0011011100110111",
									"0011011100111000",
									"0011011100111001",
									"0011011101000000",
									"0011011101000001",
									"0011011101000010",
									"0011011101000011",
									"0011011101000100",
									"0011011101000101",
									"0011011101000110",
									"0011011101000111",
									"0011011101001000",
									"0011011101001001",
									"0011011101010000",
									"0011011101010001",
									"0011011101010010",
									"0011011101010011",
									"0011011101010100",
									"0011011101010101",
									"0011011101010110",
									"0011011101010111",
									"0011011101011000",
									"0011011101011001",
									"0011011101100000",
									"0011011101100001",
									"0011011101100010",
									"0011011101100011",
									"0011011101100100",
									"0011011101100101",
									"0011011101100110",
									"0011011101100111",
									"0011011101101000",
									"0011011101101001",
									"0011011101110000",
									"0011011101110001",
									"0011011101110010",
									"0011011101110011",
									"0011011101110100",
									"0011011101110101",
									"0011011101110110",
									"0011011101110111",
									"0011011101111000",
									"0011011101111001",
									"0011011110000000",
									"0011011110000001",
									"0011011110000010",
									"0011011110000011",
									"0011011110000100",
									"0011011110000101",
									"0011011110000110",
									"0011011110000111",
									"0011011110001000",
									"0011011110001001",
									"0011011110010000",
									"0011011110010001",
									"0011011110010010",
									"0011011110010011",
									"0011011110010100",
									"0011011110010101",
									"0011011110010110",
									"0011011110010111",
									"0011011110011000",
									"0011011110011001",
									"0011100000000000",
									"0011100000000001",
									"0011100000000010",
									"0011100000000011",
									"0011100000000100",
									"0011100000000101",
									"0011100000000110",
									"0011100000000111",
									"0011100000001000",
									"0011100000001001",
									"0011100000010000",
									"0011100000010001",
									"0011100000010010",
									"0011100000010011",
									"0011100000010100",
									"0011100000010101",
									"0011100000010110",
									"0011100000010111",
									"0011100000011000",
									"0011100000011001",
									"0011100000100000",
									"0011100000100001",
									"0011100000100010",
									"0011100000100011",
									"0011100000100100",
									"0011100000100101",
									"0011100000100110",
									"0011100000100111",
									"0011100000101000",
									"0011100000101001",
									"0011100000110000",
									"0011100000110001",
									"0011100000110010",
									"0011100000110011",
									"0011100000110100",
									"0011100000110101",
									"0011100000110110",
									"0011100000110111",
									"0011100000111000",
									"0011100000111001",
									"0011100001000000",
									"0011100001000001",
									"0011100001000010",
									"0011100001000011",
									"0011100001000100",
									"0011100001000101",
									"0011100001000110",
									"0011100001000111",
									"0011100001001000",
									"0011100001001001",
									"0011100001010000",
									"0011100001010001",
									"0011100001010010",
									"0011100001010011",
									"0011100001010100",
									"0011100001010101",
									"0011100001010110",
									"0011100001010111",
									"0011100001011000",
									"0011100001011001",
									"0011100001100000",
									"0011100001100001",
									"0011100001100010",
									"0011100001100011",
									"0011100001100100",
									"0011100001100101",
									"0011100001100110",
									"0011100001100111",
									"0011100001101000",
									"0011100001101001",
									"0011100001110000",
									"0011100001110001",
									"0011100001110010",
									"0011100001110011",
									"0011100001110100",
									"0011100001110101",
									"0011100001110110",
									"0011100001110111",
									"0011100001111000",
									"0011100001111001",
									"0011100010000000",
									"0011100010000001",
									"0011100010000010",
									"0011100010000011",
									"0011100010000100",
									"0011100010000101",
									"0011100010000110",
									"0011100010000111",
									"0011100010001000",
									"0011100010001001",
									"0011100010010000",
									"0011100010010001",
									"0011100010010010",
									"0011100010010011",
									"0011100010010100",
									"0011100010010101",
									"0011100010010110",
									"0011100010010111",
									"0011100010011000",
									"0011100010011001",
									"0011100100000000",
									"0011100100000001",
									"0011100100000010",
									"0011100100000011",
									"0011100100000100",
									"0011100100000101",
									"0011100100000110",
									"0011100100000111",
									"0011100100001000",
									"0011100100001001",
									"0011100100010000",
									"0011100100010001",
									"0011100100010010",
									"0011100100010011",
									"0011100100010100",
									"0011100100010101",
									"0011100100010110",
									"0011100100010111",
									"0011100100011000",
									"0011100100011001",
									"0011100100100000",
									"0011100100100001",
									"0011100100100010",
									"0011100100100011",
									"0011100100100100",
									"0011100100100101",
									"0011100100100110",
									"0011100100100111",
									"0011100100101000",
									"0011100100101001",
									"0011100100110000",
									"0011100100110001",
									"0011100100110010",
									"0011100100110011",
									"0011100100110100",
									"0011100100110101",
									"0011100100110110",
									"0011100100110111",
									"0011100100111000",
									"0011100100111001",
									"0011100101000000",
									"0011100101000001",
									"0011100101000010",
									"0011100101000011",
									"0011100101000100",
									"0011100101000101",
									"0011100101000110",
									"0011100101000111",
									"0011100101001000",
									"0011100101001001",
									"0011100101010000",
									"0011100101010001",
									"0011100101010010",
									"0011100101010011",
									"0011100101010100",
									"0011100101010101",
									"0011100101010110",
									"0011100101010111",
									"0011100101011000",
									"0011100101011001",
									"0011100101100000",
									"0011100101100001",
									"0011100101100010",
									"0011100101100011",
									"0011100101100100",
									"0011100101100101",
									"0011100101100110",
									"0011100101100111",
									"0011100101101000",
									"0011100101101001",
									"0011100101110000",
									"0011100101110001",
									"0011100101110010",
									"0011100101110011",
									"0011100101110100",
									"0011100101110101",
									"0011100101110110",
									"0011100101110111",
									"0011100101111000",
									"0011100101111001",
									"0011100110000000",
									"0011100110000001",
									"0011100110000010",
									"0011100110000011",
									"0011100110000100",
									"0011100110000101",
									"0011100110000110",
									"0011100110000111",
									"0011100110001000",
									"0011100110001001",
									"0011100110010000",
									"0011100110010001",
									"0011100110010010",
									"0011100110010011",
									"0011100110010100",
									"0011100110010101",
									"0011100110010110",
									"0011100110010111",
									"0011100110011000",
									"0011100110011001",
									"0100000000000000",
									"0100000000000001",
									"0100000000000010",
									"0100000000000011",
									"0100000000000100",
									"0100000000000101",
									"0100000000000110",
									"0100000000000111",
									"0100000000001000",
									"0100000000001001",
									"0100000000010000",
									"0100000000010001",
									"0100000000010010",
									"0100000000010011",
									"0100000000010100",
									"0100000000010101",
									"0100000000010110",
									"0100000000010111",
									"0100000000011000",
									"0100000000011001",
									"0100000000100000",
									"0100000000100001",
									"0100000000100010",
									"0100000000100011",
									"0100000000100100",
									"0100000000100101",
									"0100000000100110",
									"0100000000100111",
									"0100000000101000",
									"0100000000101001",
									"0100000000110000",
									"0100000000110001",
									"0100000000110010",
									"0100000000110011",
									"0100000000110100",
									"0100000000110101",
									"0100000000110110",
									"0100000000110111",
									"0100000000111000",
									"0100000000111001",
									"0100000001000000",
									"0100000001000001",
									"0100000001000010",
									"0100000001000011",
									"0100000001000100",
									"0100000001000101",
									"0100000001000110",
									"0100000001000111",
									"0100000001001000",
									"0100000001001001",
									"0100000001010000",
									"0100000001010001",
									"0100000001010010",
									"0100000001010011",
									"0100000001010100",
									"0100000001010101",
									"0100000001010110",
									"0100000001010111",
									"0100000001011000",
									"0100000001011001",
									"0100000001100000",
									"0100000001100001",
									"0100000001100010",
									"0100000001100011",
									"0100000001100100",
									"0100000001100101",
									"0100000001100110",
									"0100000001100111",
									"0100000001101000",
									"0100000001101001",
									"0100000001110000",
									"0100000001110001",
									"0100000001110010",
									"0100000001110011",
									"0100000001110100",
									"0100000001110101",
									"0100000001110110",
									"0100000001110111",
									"0100000001111000",
									"0100000001111001",
									"0100000010000000",
									"0100000010000001",
									"0100000010000010",
									"0100000010000011",
									"0100000010000100",
									"0100000010000101",
									"0100000010000110",
									"0100000010000111",
									"0100000010001000",
									"0100000010001001",
									"0100000010010000",
									"0100000010010001",
									"0100000010010010",
									"0100000010010011",
									"0100000010010100",
									"0100000010010101");
  
begin

  -- Reads ROM position at every rising edge of 'clk'.
  process (clk)
  begin
	if (clk'event and clk = '1') then
  		out_rom <= memory(to_integer(unsigned(address)));
    end if;
  end process;

end architecture rom_bcd;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 2, 0, 0, 0, 2, 1, 1, 0, 1, 2, 2, 2, 0, 1, 0, 2, 1, 2, 0, 0, 0, 2, 0, -2, -2, -2, 2, 1, -2, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -2, 2, 0, 0, 1, 1, -2, -2, -2, 2, 1, 1, 0, 0, 0, -2, 1, 1, 0, -2, -2, -2, 1, -2, -2, 2, -2, -2, 2, 1, 1, 1, 0, 1, 1, -2, -2, -2, 1, 1, -2, -2, 2, 0, -2, -2, -2, 2, -2, 1, 0, -2, -2, 1, 0, 1, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, 0, 1, 2, -2, -2, -2, 1, -2, 1, 2, 1, 1, -2, -2, -2, -2, 0, 1, 0, 1, -2, -2, -2, 0, 2, -2, 1, 0, 0, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 2, 1, 1, -2, -2, 0, 0, 1, 0, 2, -2, 2, 0, -2, -2, -2, 0, 1, 1, -2, -2, 1, -2, 0, -2, -2, 0, -2, 1, 0, 0, -2, 0, 1, -2, -2, -2, -2, 1, -2, 1, 2, 0, 2, -2, 2, 0, -2, -2, 1, 1, -2, -2, -2, -2, 0, -2, -2, 0, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, 1, -2, 1, 2, 0, -2, 1, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 0, -2, -2, -2, 2, -2, 1, -2, -2, -2, 1, 0, -2, -2, -2, -2, 0, -2, -2, -2, -2, 0, -2, -2, -2, 0, -2, -2, -2, -2, 0, -2, -2, 1, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, 0, 0, -2, 2, -2, -2, -2, 0, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 0, 1, 1, 1, 2, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 1, 2, 1, 1, 0, -2, 2, 2, 0, 0, 1, 1, 1, 2, 1, 2, 0, 0, 2, 2, 0, -2, 1, 1, 1, 1, 1, 2, 1, 0, 1, 0, 1, 2, 2, -2, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, -2, -2, -2, -2, 1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 0, 2, 2, 1, 0, 0, -2, 0, -2, 1, 1, 0, -2, -2, 2, 0, 1, 1, -2, 2, 0, 0, 0, -2, 2, -2, 1, 2, 0, 0, 1, 1, 0, 2, 0, 1, -2, -2, 1, 1, 1, 2, -2, 0, 1, 0, -2, -2, 0, 1, 0, 2, 2, 1, 0, 2, 2, -2, 0, 1, -2, -2, 1, 1, 1, 2, 1, -2, 2, 2, 1, 0, -2, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, 0, -2, -2, 0, -2, -2, -2, -2, -2, 2, 1, 1, 1, -2, -2, -2, -2, 0, 0, -2, -2, -2, 1, -2, -2, -2, 2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 2, -2, -2, -2, 0, -2, -2, 1, 1, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, 1, 2, 1, -2, 2, 1, -2, -2, -2, -2, -2, -2, -2, 1, 0, -2, -2, -2, 0, 2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, 2, -2, -2, 1, 0, 1, 2, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, 2, 0, -2, 0, -2, -2, -2, -2, -2, -2, 1, -2, 0, -2, -2, -2, -2, 0, 1, 1, 1, -2, -2, -2, -2, 2, -2, -2, 0, -2, -2, -2, 2, -2, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, 0, -2, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 1, 1, -2, -2, -2, -2, 1, 2, 0, -2, 0, -2, -2, -2, 0, -2, -2, -2, -2, 1, -2, -2, -2, 2, -2, -2, -2, 2, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, 0, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, 1, -2, -2, 0, -2, -2, -2, -2, -2, 1, -2, -2, 2, 1, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((1068534, 53900, 1921424, 281086, 791101, 21938, 41380, 84674, 2370806, 74627, 4285, 96825, 1397682, 75658, 29734, 61504, 73568, 3502, 88251, 7032, 117678, 94858, 105794, 372672, 486055, 4285, 614654, 1546709, 1843567, 1384693, 2929, 5238, 102266, 1838506, 1666785, 63352, 65871, 899818, 975816, 69570, 3502, 1396319, 1220432, 2929, 1521762, 1476057, 1675628, 5238, 118152, 97702, 2743984, 94273, 3502, 2929, 4285, 608518, 68006, 530958, 3502, 56223, 4285, 167894, 255505, 140595, 4285, 20361, -8192, -8192, -8192, 4285, 92000, -8192, 901721, 100591, 106756, 2088300, 2335336, 1565589, 1512705, 79305, 83404, 13251, 21666, 11893, 4285, 4285, 2929, 48313, 493459, 534851, 611976, 103572, 2203237, 1219468, 1360628, -8192, 5238, 482561, 424355, 45777, 50504, -8192, -8192, -8192, 3502, 85565, 93988, 962686, 1020360, 1188529, -8192, 86782, 92411, 349288, -8192, -8192, -8192, 59043, -8192, -8192, 2929, -8192, -8192, 2929, 81759, 78865, 82338, 1765031, 91312, 28485, -8192, -8192, -8192, 91175, 95666, -8192, -8192, 5238, 895732, -8192, -8192, -8192, 4285, -8192, 58176, 212596, -8192, -8192, 78140, 1207186, 80773, -8192, -8192, -8192, -8192, 740171, -8192, -8192, -8192, -8192, -8192, 943467, 68889, 2929, -8192, -8192, -8192, 33790, -8192, 32570, 4285, 37287, 39364, -8192, -8192, -8192, -8192, 1718608, 101937, 1888563, 105102, -8192, -8192, -8192, 902499, 4285, -8192, 67479, 853722, 321639, -8192, -8192, -8192, -8192, -8192, 107665, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 18389, -8192, -8192, -8192, -8192, -8192, 4285, 83525, 78188, -8192, -8192, 1136292, 655669, 70105, 610515, 4285, -8192, 5238, 704904, -8192, -8192, -8192, 2259425, 102097, 99729, -8192, -8192, 57449, -8192, 82110, -8192, -8192, 2051331, -8192, 111637, 2096244, 1987557, -8192, 245826, 37578, -8192, -8192, -8192, -8192, 108245, -8192, 104595, 2929, 2636691, 3502, -8192, 2929, 2071333, -8192, -8192, 95475, 56006, -8192, -8192, -8192, -8192, 142783, -8192, -8192, 773133, -8192, 50822, -8192, -8192, -8192, -8192, 110155, -8192, -8192, -8192, -8192, -8192, -8192, 41870, -8192, 66952, 2929, 1228700, -8192, 70916, 1348899, 71559, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 1738884, -8192, -8192, 24237, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 99796, -8192, -8192, 5238, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 5238, -8192, -8192, -8192, 82899, -8192, -8192, -8192, -8192, -8192, 332448, -8192, -8192, -8192, 3502, -8192, 104079, -8192, -8192, -8192, 104844, 2422900, -8192, -8192, -8192, -8192, 1391100, -8192, -8192, -8192, -8192, 2089431, -8192, -8192, -8192, 2476024, -8192, -8192, -8192, -8192, 947673, -8192, -8192, 103373, -8192, -8192, -8192, 672516, -8192, -8192, -8192, 101704, -8192, -8192, -8192, -8192, -8192, -8192, 33623, -8192, -8192, -8192, 83638, -8192, -8192, 681558, 779853, -8192, 4285, -8192, -8192, -8192, 780466, -8192, -8192, 91826, -8192, -8192, -8192, -8192, 66986, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192),
                (1396964, 52445, 2136951, 360793, 873318, 22101, 494865, 90605, 2576813, 81727, 4285, 99480, 1680810, 62390, 75233, 68550, 4285, 88865, 283114, 8402, 141734, 41507, 574439, 37458, 5238, 79942, 91924, 1034991, 1344172, 62960, 4285, 82454, 88258, 1069856, -8192, 3502, 3502, 1873052, 1630963, 102629, 116699, 101353, 5238, 77526, 2929, 1906788, 1608546, 3502, 2929, 1592565, -8192, 28401, 34148, 31894, 39975, 93355, 2929, 107533, 1429727, 104680, 2786968, 100009, 3502, 2929, -8192, 1249558, 1157240, 614799, 695921, 499989, 4285, 3502, 60512, 93687, 1680577, 77228, 5238, 37744, 79771, 21345, 7062, 2500786, 2336452, 93922, 97721, 109654, 110798, 456056, 373773, 830407, 718956, 56607, 60032, -8192, -8192, -8192, -8192, 102324, 1923405, 1722570, 108117, 105352, 2043439, 1199082, 99745, 95333, 5238, 184353, 276385, 154548, 2929, 3502, 83526, 1315635, 1073018, -8192, 1192560, -8192, 115136, 85677, 1153443, -8192, -8192, 3502, 1661947, 87455, 89903, -8192, 2929, 1110345, 921600, 1053861, -8192, 3502, -8192, 99106, 2929, 2363879, 2212355, 17318, 19997, 102400, 4285, 1480062, 96544, -8192, -8192, 101198, 101599, 33462, 2929, -8192, 372575, 86384, 1543915, -8192, -8192, 365855, 49452, 451599, 5238, 4285, 57494, 285704, 3502, 2929, -8192, 734150, 56755, -8192, -8192, 46982, 49621, 43732, 4285, 48220, -8192, 4285, 5238, 36213, 291329, -8192, -8192, -8192, -8192, -8192, 103873, -8192, -8192, -8192, 83513, -8192, 1858864, -8192, -8192, 1579471, -8192, -8192, -8192, -8192, -8192, 4285, 44317, 42925, 46145, -8192, -8192, -8192, -8192, 2394349, 2428555, -8192, -8192, -8192, 55846, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, -8192, 61804, -8192, -8192, -8192, 4285, -8192, -8192, -8192, 1814588, -8192, -8192, 94790, 97731, -8192, -8192, -8192, 105749, -8192, -8192, -8192, 71148, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 60561, -8192, -8192, -8192, -8192, 1643401, -8192, -8192, -8192, -8192, -8192, -8192, 71492, 4285, 76065, -8192, 5238, 67374, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 107395, 2293642, -8192, -8192, -8192, 734596, 5238, -8192, -8192, -8192, -8192, -8192, 1766896, -8192, -8192, -8192, 535669, -8192, -8192, -8192, -8192, -8192, 75813, 2929, -8192, -8192, 109570, 2887680, 107801, 2929, 112843, -8192, 110124, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 610864, 2929, 756591, -8192, 650576, -8192, -8192, -8192, -8192, -8192, -8192, 33712, -8192, 365427, -8192, -8192, -8192, -8192, 1349285, 86349, 83268, 82330, -8192, -8192, -8192, -8192, 5238, -8192, -8192, 738533, -8192, -8192, -8192, 2929, -8192, -8192, -8192, 112269, -8192, -8192, -8192, -8192, 107039, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 3502, -8192, -8192, -8192, -8192, 2049003, -8192, 1998858, 2929, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 14840, -8192, -8192, -8192, -8192, 29225, 34143, -8192, -8192, -8192, -8192, 74774, 2929, 1555822, -8192, 1479106, -8192, -8192, -8192, 2204838, -8192, -8192, -8192, -8192, 46115, -8192, -8192, -8192, 5238, -8192, -8192, -8192, 5238, -8192, 57977, -8192, -8192, -8192, 43748, -8192, -8192, -8192, -8192, 1644435, -8192, -8192, -8192, 92944, 2267366, -8192, -8192, -8192, -8192, -8192, 20111, -8192, -8192, 226903, -8192, -8192, -8192, -8192, -8192, 110675, -8192, -8192, 2929, 113390, -8192, -8192, -8192, 610092, -8192, -8192, -8192, 86275, -8192, -8192, -8192, -8192, 74849, -8192, -8192, -8192, 93043, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192),
                (2084370, 53338, 2887680, 536081, 1187550, -8192, -8192, -8192, -8192, 99886, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((1226, 561, 1329, 1049, 126, 449, 1270, 1107, 1359, 1336, 475, 200, 914, 942, 112, 39, 390, 1004, 102, 225, 1232, 485, 1180, 1350, 1008, 203, 1270, 474, 32, 129, 890, 1097, 179, 222, 1212, 637, 1258, 1142, 195, 1361, 1133, 863, 1322, 244, 1214, 1345, 822, 428, 1300, 1289, 1364, 1361, 898, 327, 1317, 234, 11, 47, 863, 178, 1214, 390, 16, 35, 1066, 759, 0, 0, 1365, 297, 4, 0, 738, 82, 569, 941, 140, 91, 910, 352, 1016, 871, 1327, 1317, 216, 1011, 1342, 730, 1329, 1092, 228, 427, 1224, 488, 17, 0, 759, 37, 465, 228, 1241, 248, 1109, 0, 359, 137, 883, 1264, 597, 837, 1365, 341, 1150, 745, 0, 0, 1365, 759, 1365, 1365, 152, 1155, 0, 893, 1328, 455, 1268, 44, 683, 780, 1365, 1092, 0, 926, 1343, 1274, 525, 735, 76, 455, 1252, 0, 341, 0, 993, 964, 0, 0, 455, 840, 161, 228, 1365, 228, 1170, 796, 1365, 273, 1138, 683, 1365, 37, 503, 869, 0, 607, 0, 1247, 1365, 1358, 640, 273, 1252, 1138, 228, 607, 1365, 10, 254, 956, 41, 455, 1365, 1365, 1121, 710, 1365, 114, 1260, 683, 0, 0, 1092, 819, 0, 76, 910, 1365, 683, 1365, 546, 683, 0, 1342, 683, 1365, 546, 91, 910, 1144, 1358, 621, 1365, 1365, 195, 79, 2, 13, 423, 0, 1109, 683, 1365, 0, 1365, 341, 20, 114, 1024, 683, 72, 0, 512, 0, 819, 1223, 1365, 931, 1341, 1205, 0, 4, 228, 819, 0, 1024, 1365, 1345, 1365, 1363, 1090, 98, 1341, 1365, 1267, 853, 1365, 0, 1241, 585, 1092, 1024, 0, 1365, 1187, 341, 1365, 1250, 1365, 910, 1365, 1365, 228, 0, 303, 910, 0, 1365, 910, 1062, 1365, 19, 455, 1365, 1312, 1062, 1365, 341, 1268, 910, 1365, 1365, 455, 683, 0, 0, 455, 0, 273, 1330, 910, 0, 210, 910, 0, 455, 41, 1365, 910, 455, 0, 910, 1365, 1365, 910, 1237, 1365, 1365, 993, 341, 1365, 341, 0, 1024, 1365, 0, 455, 303, 0, 1365, 1062, 455, 0, 1365, 1024, 1365, 1024, 0, 341, 0, 124, 0, 910, 1365, 1222, 1092, 1365, 1365, 1138, 1365, 1170, 910, 1365, 0, 62, 0, 228, 683, 0, 1365, 1311, 683, 1365, 455, 910, 0, 171, 455, 0, 0, 195, 1195, 1365, 1365, 910, 1271, 1365, 819, 1365, 0, 171, 455, 0, 171, 0, 0, 455, 195, 0, 0, 455, 124, 0, 0, 455, 1252, 1365, 0, 72, 455, 0, 1365, 1297, 910, 1365, 33, 1, 0, 273, 0, 910, 0, 49, 455, 0, 23, 0, 0, 455, 1365, 1353, 910, 1365, 0, 0, 0, 0, 1365, 1365, 0, 0, 0, 0, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 910, 910, 1365, 1365, 546, 546, 683, 683, 1365, 1365, 546, 546, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 1024, 1024, 683, 683, 0, 0, 1365, 1365, 0, 0, 819, 819, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1092, 1092, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 910, 910, 0, 0, 1365, 1365, 910, 910, 455, 455, 1365, 1365, 1365, 1365, 683, 683, 0, 0, 910, 910, 0, 0, 910, 910, 0, 0, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 1365, 1365, 341, 341, 0, 0, 1024, 1024, 1365, 1365, 0, 0, 0, 0, 910, 910, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 455, 455, 910, 910, 0, 0, 1365, 1365, 1365, 1365, 819, 819, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 455, 455, 0, 0, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 0, 0, 910, 910, 0, 0, 455, 455, 0, 0, 0, 0, 0, 0, 455, 455, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 819, 819, 819, 819, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365),
                (1091, 403, 1322, 932, 134, 318, 1290, 1063, 1358, 1331, 433, 181, 1094, 29, 368, 1098, 144, 780, 105, 178, 1292, 968, 1349, 1308, 208, 31, 344, 908, 83, 1282, 765, 398, 1226, 523, 1365, 435, 74, 251, 970, 812, 1343, 1344, 460, 1363, 1080, 443, 1270, 88, 864, 182, 1365, 47, 394, 1153, 104, 60, 661, 139, 945, 1278, 1364, 1353, 744, 241, 1365, 431, 1265, 149, 8, 36, 564, 275, 1280, 420, 1302, 993, 168, 495, 20, 65, 1163, 30, 575, 332, 1112, 188, 975, 96, 834, 127, 662, 91, 1138, 878, 0, 114, 975, 12, 226, 73, 826, 1289, 410, 41, 410, 1229, 205, 225, 6, 22, 1083, 226, 8, 48, 645, 0, 1161, 0, 1084, 1350, 910, 293, 1303, 1052, 1358, 556, 1336, 1365, 1121, 661, 1276, 152, 1365, 683, 1365, 1364, 1133, 534, 1344, 1024, 1358, 1325, 293, 1024, 152, 1365, 512, 124, 910, 1348, 975, 0, 1241, 853, 124, 0, 819, 228, 1138, 5, 208, 69, 1050, 1323, 735, 195, 1365, 55, 569, 1365, 0, 1228, 1360, 1320, 455, 195, 1365, 352, 16, 62, 1062, 1365, 683, 1183, 341, 1365, 455, 228, 1138, 0, 405, 1365, 186, 1365, 546, 431, 0, 182, 1365, 0, 416, 18, 372, 1138, 85, 0, 819, 455, 1365, 1260, 728, 228, 1062, 0, 420, 1092, 0, 1365, 1040, 0, 1365, 621, 1365, 1365, 819, 0, 1365, 546, 1195, 0, 410, 1365, 956, 341, 1365, 5, 147, 520, 51, 0, 210, 607, 0, 0, 341, 780, 0, 0, 546, 1365, 683, 76, 683, 1365, 780, 341, 1365, 0, 546, 910, 1365, 1365, 455, 683, 1365, 0, 38, 247, 7, 0, 956, 683, 1365, 993, 195, 910, 1365, 683, 1365, 455, 68, 228, 910, 1365, 1073, 780, 1365, 0, 1365, 1073, 1365, 149, 0, 85, 585, 455, 0, 910, 0, 1024, 1365, 18, 303, 0, 683, 1341, 1365, 1363, 951, 144, 1365, 390, 0, 0, 683, 1365, 910, 910, 1365, 910, 1365, 1365, 1293, 975, 1365, 195, 1365, 455, 0, 455, 0, 1365, 1229, 455, 1315, 910, 1365, 0, 455, 74, 1, 16, 910, 455, 1365, 0, 455, 88, 0, 0, 607, 0, 1365, 1365, 1222, 683, 1365, 0, 171, 0, 341, 0, 146, 303, 0, 0, 455, 455, 0, 0, 455, 0, 144, 0, 273, 0, 273, 70, 0, 19, 683, 0, 1365, 0, 273, 0, 455, 1365, 910, 341, 0, 1365, 1024, 0, 119, 546, 0, 1365, 1092, 2, 101, 910, 0, 1092, 1365, 1365, 1325, 1163, 1365, 455, 1365, 137, 0, 1229, 1365, 1365, 910, 0, 124, 455, 0, 1365, 1241, 910, 1365, 0, 54, 0, 341, 910, 0, 0, 91, 455, 0, 137, 0, 1289, 1365, 1365, 910, 1365, 1297, 910, 1365, 1365, 1285, 1365, 1297, 910, 1365, 49, 0, 0, 455, 36, 0, 1357, 1365, 1365, 1208, 910, 1365, 1092, 683, 1343, 1365, 1365, 910, 18, 0, 0, 455, 1365, 1351, 910, 1365, 1365, 1351, 910, 1365, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 0, 0, 819, 819, 455, 455, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 546, 546, 1365, 1365, 341, 341, 1365, 1365, 0, 0, 0, 0, 0, 0, 546, 546, 1365, 1365, 683, 683, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 0, 0, 0, 0, 683, 683, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 910, 910, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 455, 455, 0, 0, 0, 0, 1365, 1365, 683, 683, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 455, 455, 341, 341, 0, 0, 0, 0, 546, 546, 0, 0, 910, 910, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 910, 910, 0, 0, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1092, 1092, 683, 683, 1365, 1365, 1365, 1365, 910, 910, 0, 0, 1365, 1365, 910, 910, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 455, 455, 455, 455, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 341, 341, 341, 341, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365),
                (682, 204, 1329, 617, 85, 168, 1328, 20, 301, 1131, 1365, 1354, 520, 168, 168, 1328, 1328, 20, 20, 301, 301, 1365, 1365, 1354, 1354, 520, 520, 168, 168, 168, 168, 1328, 1328, 1328, 1328, 20, 20, 20, 20, 301, 301, 301, 301, 1365, 1365, 1365, 1365, 1354, 1354, 1354, 1354, 520, 520, 520, 520, 168, 168, 168, 168, 168, 168, 168, 168, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 20, 20, 20, 20, 20, 20, 20, 20, 301, 301, 301, 301, 301, 301, 301, 301, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 520, 520, 520, 520, 520, 520, 520, 520, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 1328, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 301, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 1354, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 520, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 7, 5, 15, 13, 23, 9, 49, 39, 11, 27, 21, 19, 61, 55, 17, 35, 69, 65, 81, 31, 45, 167, 25, 97, 85, 29, 177, 103, 33, 109, 93, 127, 133, 37, 183, 117, 161, 283, 41, 43, 209, 147, 123, 315, 47, 77, 299, 51, 247, 253, 53, 73, 235, 57, 215, 141, 59, 229, 155, 63, 241, 301, 129, 67, 423, 425, 427, 71, 415, 429, 79, 225, 75, 91, 195, 297, 139, 137, 107, 83, 203, 277, 231, 87, 267, 89, 323, 159, 207, 201, 245, 95, 365, 431, 101, 281, 99, 113, 313, -1, -1, 433, 105, 165, 121, 279, 157, 111, 435, 193, 197, 115, 437, -1, -1, 119, 439, 441, 325, -1, -1, 125, 343, 131, 333, 369, 173, 145, 443, -1, -1, 135, 347, -1, -1, 153, 295, -1, -1, 445, 143, 447, 199, 175, 449, 451, 149, 151, 327, -1, -1, -1, -1, 259, 453, -1, -1, -1, -1, 379, 163, 181, 455, -1, -1, 169, 457, 349, 171, 189, 307, -1, -1, -1, -1, 353, 179, 205, 383, -1, -1, 459, 185, 187, 461, 309, 335, 191, 463, -1, -1, -1, -1, 305, 465, -1, -1, 467, 469, -1, -1, 263, 471, 473, 475, -1, -1, 211, 401, 213, 477, 479, 331, 217, 405, 339, 219, 481, 221, 223, 483, -1, -1, 227, 391, 337, 485, 487, 387, 489, 233, -1, -1, 237, 491, 239, 371, 329, 493, 397, 243, 495, 497, -1, -1, 249, 499, 359, 251, 273, 375, 501, 255, 257, 503, 505, 311, 261, 507, -1, -1, 509, 265, -1, -1, 269, 511, 271, 513, -1, -1, 515, 275, 517, 519, 521, 523, -1, -1, 321, 525, 419, 285, 287, 527, 293, 289, 291, 529, -1, -1, 531, 533, -1, -1, -1, -1, 395, 535, 537, 303, 539, 541, -1, -1, 543, 545, -1, -1, 547, 549, 551, 553, 317, 555, 557, 319, -1, -1, 559, 561, 563, 565, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 567, 341, 569, 571, 573, 345, -1, -1, -1, -1, 575, 351, 577, 579, 581, 355, 583, 357, -1, -1, 585, 361, 363, 587, 589, 591, 593, 367, -1, -1, -1, -1, 373, 595, -1, -1, 377, 597, 599, 601, 603, 381, -1, -1, 385, 605, -1, -1, 389, 607, -1, -1, 393, 609, -1, -1, -1, -1, 611, 399, 613, 615, 617, 403, 619, 621, 407, 411, 623, 409, 625, 627, 629, 413, 631, 633, 417, 635, 637, 639, 641, 421, 643, 645, 647, 649, 651, 653, 655, 657, 659, 661, -1, -1, 663, 665, 667, 669, -1, -1, 671, 673, -1, -1, 675, 677, 679, 681, 683, 685, -1, -1, 687, 689, 691, 693, -1, -1, 695, 697, 699, 701, 703, 705, -1, -1, -1, -1, -1, -1, -1, -1, 707, 709, -1, -1, -1, -1, 711, 713, -1, -1, 715, 717, -1, -1, -1, -1, 719, 721, -1, -1, 723, 725, -1, -1, 727, 729, 731, 733, 735, 737, 739, 741, 743, 745, 747, 749, -1, -1, -1, -1, 751, 753, -1, -1, 755, 757, -1, -1, -1, -1, -1, -1, -1, -1, 759, 761, 763, 765, -1, -1, -1, -1, -1, -1, -1, -1, 767, 769, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 771, 773, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 775, 777, -1, -1, -1, -1, -1, -1, 779, 781, -1, -1, -1, -1, 783, 785, -1, -1, 787, 789, 791, 793, -1, -1, -1, -1, -1, -1, -1, -1, 795, 797, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 799, 801, -1, -1, -1, -1, 803, 805, -1, -1, -1, -1, 807, 809, -1, -1, -1, -1, 811, 813, -1, -1, -1, -1, 815, 817, 819, 821, 823, 825, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, -1, -1, -1, -1, -1, -1, -1, -1, 847, 849, 851, 853, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 855, 857, 859, 861, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 863, 865, 867, 869, 871, 873, 875, 877, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 879, 881, 883, 885, -1, -1, -1, -1, -1, -1, -1, -1, 887, 889, 891, 893, 895, 897, 899, 901, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, 951, 953, 955, 957, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 959, 961, 963, 965, 967, 969, 971, 973, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 13, 17, 21, 9, 59, 43, 11, 35, 39, 67, 15, 29, 25, 19, 51, 77, 139, 23, 171, 149, 87, 111, 27, 31, 103, 127, 33, 75, 119, 47, 485, 37, 97, 55, 73, 41, 231, 421, 57, 405, 45, 49, 123, 243, 65, 189, 487, 107, 53, 163, 177, 291, 83, 195, 117, 61, 305, 135, 63, 81, 489, 95, 289, 69, 265, 159, 71, 89, 283, 143, 259, 181, 199, 79, 393, 247, 223, 357, 85, 93, 145, 279, 209, 201, 157, 167, 91, 329, 193, -1, -1, -1, -1, 377, 99, 239, 101, 397, 155, 235, 105, 391, 229, 109, 399, 371, 227, 113, 339, 301, 115, 491, 275, 493, 183, 445, 121, -1, -1, 125, 437, 153, 315, 495, 129, 131, 133, 257, 497, 187, 499, 441, 137, 147, 413, 141, 447, 317, 205, 277, 375, -1, -1, 389, 185, 331, 151, 501, 207, 221, 337, -1, -1, 385, 249, 425, 161, 213, 253, 319, 165, 369, 503, 361, 169, -1, -1, 173, 321, 217, 175, 295, 505, 179, 431, 435, 263, -1, -1, -1, -1, 507, 483, -1, -1, 509, 191, 511, 251, -1, -1, 197, 513, -1, -1, -1, -1, 417, 203, 387, 327, 515, 517, 519, 521, 403, 211, -1, -1, 523, 215, -1, -1, 525, 219, 527, 529, -1, -1, 531, 225, -1, -1, 533, 299, -1, -1, 535, 233, 537, 539, 455, 237, -1, -1, 541, 241, -1, -1, 543, 245, -1, -1, 545, 547, 549, 551, -1, -1, 553, 255, -1, -1, -1, -1, 261, 555, -1, -1, -1, -1, 557, 267, 269, 347, 559, 271, 273, 561, -1, -1, -1, -1, -1, -1, 281, 359, -1, -1, 563, 285, 287, 565, -1, -1, -1, -1, 293, 567, -1, -1, 297, 569, -1, -1, -1, -1, 411, 303, -1, -1, 307, 457, 353, 309, 311, 571, 313, 573, 575, 577, 579, 581, 583, 585, 587, 589, 465, 323, 325, 591, 367, 593, -1, -1, -1, -1, 595, 333, 597, 335, -1, -1, -1, -1, 341, 469, 345, 343, -1, -1, -1, -1, 349, 599, 601, 351, -1, -1, 603, 355, 605, 607, 609, 363, -1, -1, -1, -1, 365, 611, -1, -1, -1, -1, -1, -1, 613, 373, -1, -1, -1, -1, 379, 615, 383, 381, -1, -1, -1, -1, 617, 619, -1, -1, 621, 623, -1, -1, 625, 395, 627, 629, -1, -1, 451, 401, 631, 633, -1, -1, 473, 407, 409, 635, 481, 637, -1, -1, 415, 639, 641, 643, 645, 419, -1, -1, 647, 423, 649, 651, 653, 427, 655, 429, -1, -1, 657, 433, -1, -1, -1, -1, 439, 659, 661, 663, 477, 443, 665, 667, -1, -1, 669, 449, 671, 673, 453, 675, -1, -1, -1, -1, 459, 677, 679, 461, 463, 681, 683, 685, 467, 687, 689, 691, 471, 693, -1, -1, 695, 475, 697, 699, 701, 479, 703, 705, 707, 709, -1, -1, 711, 713, 715, 717, 719, 721, -1, -1, -1, -1, 723, 725, -1, -1, -1, -1, 727, 729, -1, -1, 731, 733, -1, -1, 735, 737, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 739, 741, -1, -1, -1, -1, -1, -1, -1, -1, 743, 745, 747, 749, 751, 753, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 755, 757, 759, 761, -1, -1, 763, 765, -1, -1, -1, -1, -1, -1, 767, 769, 771, 773, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 775, 777, -1, -1, 779, 781, -1, -1, 783, 785, -1, -1, 787, 789, 791, 793, 795, 797, 799, 801, -1, -1, -1, -1, 803, 805, -1, -1, -1, -1, -1, -1, -1, -1, 807, 809, -1, -1, -1, -1, -1, -1, -1, -1, 811, 813, 815, 817, 819, 821, -1, -1, -1, -1, -1, -1, 823, 825, -1, -1, -1, -1, 827, 829, -1, -1, -1, -1, 831, 833, -1, -1, -1, -1, 835, 837, 839, 841, 843, 845, -1, -1, -1, -1, -1, -1, 847, 849, 851, 853, 855, 857, -1, -1, -1, -1, 859, 861, -1, -1, -1, -1, -1, -1, 863, 865, 867, 869, 871, 873, 875, 877, -1, -1, -1, -1, -1, -1, -1, -1, 879, 881, 883, 885, 887, 889, 891, 893, 895, 897, 899, 901, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 951, 953, 955, 957, 959, 961, 963, 965, -1, -1, -1, -1, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, 13, 15, 17, 19, 11, 21, 23, 25, 27, 29, 31, 33, 35, 37, 39, 41, 43, 45, 47, 49, 51, 53, 55, 57, 59, 61, 63, 65, 67, 69, 71, 73, 75, 77, 79, 81, 83, 85, 87, 89, 91, 93, 95, 97, 99, 101, 103, 105, 107, 109, 111, 113, 115, 117, 119, 121, 123, 125, 127, 129, 131, 133, 135, 137, 139, 141, 143, 145, 147, 149, 151, 153, 155, 157, 159, 161, 163, 165, 167, 169, 171, 173, 175, 177, 179, 181, 183, 185, 187, 189, 191, 193, 195, 197, 199, 201, 203, 205, 207, 209, 211, 213, 215, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 237, 239, 241, 243, 245, 247, 249, 251, 253, 255, 257, 259, 261, 263, 265, 267, 269, 271, 273, 275, 277, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 341, 343, 345, 347, 349, 351, 353, 355, 357, 359, 361, 363, 365, 367, 369, 371, 373, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 415, 417, 419, 421, 423, 425, 427, 429, 431, 433, 435, 437, 439, 441, 443, 445, 447, 449, 451, 453, 455, 457, 459, 461, 463, 465, 467, 469, 471, 473, 475, 477, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, 511, 513, 515, 517, 519, 521, 523, 525, 527, 529, 531, 533, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 555, 557, 559, 561, 563, 565, 567, 569, 571, 573, 575, 577, 579, 581, 583, 585, 587, 589, 591, 593, 595, 597, 599, 601, 603, 605, 607, 609, 611, 613, 615, 617, 619, 621, 623, 625, 627, 629, 631, 633, 635, 637, 639, 641, 643, 645, 647, 649, 651, 653, 655, 657, 659, 661, 663, 665, 667, 669, 671, 673, 675, 677, 679, 681, 683, 685, 687, 689, 691, 693, 695, 697, 699, 701, 703, 705, 707, 709, 711, 713, 715, 717, 719, 721, 723, 725, 727, 729, 731, 733, 735, 737, 739, 741, 743, 745, 747, 749, 751, 753, 755, 757, 759, 761, 763, 765, 767, 769, 771, 773, 775, 777, 779, 781, 783, 785, 787, 789, 791, 793, 795, 797, 799, 801, 803, 805, 807, 809, 811, 813, 815, 817, 819, 821, 823, 825, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, 847, 849, 851, 853, 855, 857, 859, 861, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, 887, 889, 891, 893, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 895, 897, 899, 901, 903, 905, 907, 909, 911, 913, 915, 917, 919, 921, 923, 925, 927, 929, 931, 933, 935, 937, 939, 941, 943, 945, 947, 949, 951, 953, 955, 957, 959, 961, 963, 965, 967, 969, 971, 973, 975, 977, 979, 981, 983, 985, 987, 989, 991, 993, 995, 997, 999, 1001, 1003, 1005, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 8, 6, 16, 14, 24, 10, 50, 40, 12, 28, 22, 20, 62, 56, 18, 36, 70, 66, 82, 32, 46, 168, 26, 98, 86, 30, 178, 104, 34, 110, 94, 128, 134, 38, 184, 118, 162, 284, 42, 44, 210, 148, 124, 316, 48, 78, 300, 52, 248, 254, 54, 74, 236, 58, 216, 142, 60, 230, 156, 64, 242, 302, 130, 68, 424, 426, 428, 72, 416, 430, 80, 226, 76, 92, 196, 298, 140, 138, 108, 84, 204, 278, 232, 88, 268, 90, 324, 160, 208, 202, 246, 96, 366, 432, 102, 282, 100, 114, 314, -1, -1, 434, 106, 166, 122, 280, 158, 112, 436, 194, 198, 116, 438, -1, -1, 120, 440, 442, 326, -1, -1, 126, 344, 132, 334, 370, 174, 146, 444, -1, -1, 136, 348, -1, -1, 154, 296, -1, -1, 446, 144, 448, 200, 176, 450, 452, 150, 152, 328, -1, -1, -1, -1, 260, 454, -1, -1, -1, -1, 380, 164, 182, 456, -1, -1, 170, 458, 350, 172, 190, 308, -1, -1, -1, -1, 354, 180, 206, 384, -1, -1, 460, 186, 188, 462, 310, 336, 192, 464, -1, -1, -1, -1, 306, 466, -1, -1, 468, 470, -1, -1, 264, 472, 474, 476, -1, -1, 212, 402, 214, 478, 480, 332, 218, 406, 340, 220, 482, 222, 224, 484, -1, -1, 228, 392, 338, 486, 488, 388, 490, 234, -1, -1, 238, 492, 240, 372, 330, 494, 398, 244, 496, 498, -1, -1, 250, 500, 360, 252, 274, 376, 502, 256, 258, 504, 506, 312, 262, 508, -1, -1, 510, 266, -1, -1, 270, 512, 272, 514, -1, -1, 516, 276, 518, 520, 522, 524, -1, -1, 322, 526, 420, 286, 288, 528, 294, 290, 292, 530, -1, -1, 532, 534, -1, -1, -1, -1, 396, 536, 538, 304, 540, 542, -1, -1, 544, 546, -1, -1, 548, 550, 552, 554, 318, 556, 558, 320, -1, -1, 560, 562, 564, 566, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 568, 342, 570, 572, 574, 346, -1, -1, -1, -1, 576, 352, 578, 580, 582, 356, 584, 358, -1, -1, 586, 362, 364, 588, 590, 592, 594, 368, -1, -1, -1, -1, 374, 596, -1, -1, 378, 598, 600, 602, 604, 382, -1, -1, 386, 606, -1, -1, 390, 608, -1, -1, 394, 610, -1, -1, -1, -1, 612, 400, 614, 616, 618, 404, 620, 622, 408, 412, 624, 410, 626, 628, 630, 414, 632, 634, 418, 636, 638, 640, 642, 422, 644, 646, 648, 650, 652, 654, 656, 658, 660, 662, -1, -1, 664, 666, 668, 670, -1, -1, 672, 674, -1, -1, 676, 678, 680, 682, 684, 686, -1, -1, 688, 690, 692, 694, -1, -1, 696, 698, 700, 702, 704, 706, -1, -1, -1, -1, -1, -1, -1, -1, 708, 710, -1, -1, -1, -1, 712, 714, -1, -1, 716, 718, -1, -1, -1, -1, 720, 722, -1, -1, 724, 726, -1, -1, 728, 730, 732, 734, 736, 738, 740, 742, 744, 746, 748, 750, -1, -1, -1, -1, 752, 754, -1, -1, 756, 758, -1, -1, -1, -1, -1, -1, -1, -1, 760, 762, 764, 766, -1, -1, -1, -1, -1, -1, -1, -1, 768, 770, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 772, 774, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 776, 778, -1, -1, -1, -1, -1, -1, 780, 782, -1, -1, -1, -1, 784, 786, -1, -1, 788, 790, 792, 794, -1, -1, -1, -1, -1, -1, -1, -1, 796, 798, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 800, 802, -1, -1, -1, -1, 804, 806, -1, -1, -1, -1, 808, 810, -1, -1, -1, -1, 812, 814, -1, -1, -1, -1, 816, 818, 820, 822, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, -1, -1, -1, -1, -1, -1, -1, -1, 848, 850, 852, 854, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 856, 858, 860, 862, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 864, 866, 868, 870, 872, 874, 876, 878, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 880, 882, 884, 886, -1, -1, -1, -1, -1, -1, -1, -1, 888, 890, 892, 894, 896, 898, 900, 902, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, 952, 954, 956, 958, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 960, 962, 964, 966, 968, 970, 972, 974, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 14, 18, 22, 10, 60, 44, 12, 36, 40, 68, 16, 30, 26, 20, 52, 78, 140, 24, 172, 150, 88, 112, 28, 32, 104, 128, 34, 76, 120, 48, 486, 38, 98, 56, 74, 42, 232, 422, 58, 406, 46, 50, 124, 244, 66, 190, 488, 108, 54, 164, 178, 292, 84, 196, 118, 62, 306, 136, 64, 82, 490, 96, 290, 70, 266, 160, 72, 90, 284, 144, 260, 182, 200, 80, 394, 248, 224, 358, 86, 94, 146, 280, 210, 202, 158, 168, 92, 330, 194, -1, -1, -1, -1, 378, 100, 240, 102, 398, 156, 236, 106, 392, 230, 110, 400, 372, 228, 114, 340, 302, 116, 492, 276, 494, 184, 446, 122, -1, -1, 126, 438, 154, 316, 496, 130, 132, 134, 258, 498, 188, 500, 442, 138, 148, 414, 142, 448, 318, 206, 278, 376, -1, -1, 390, 186, 332, 152, 502, 208, 222, 338, -1, -1, 386, 250, 426, 162, 214, 254, 320, 166, 370, 504, 362, 170, -1, -1, 174, 322, 218, 176, 296, 506, 180, 432, 436, 264, -1, -1, -1, -1, 508, 484, -1, -1, 510, 192, 512, 252, -1, -1, 198, 514, -1, -1, -1, -1, 418, 204, 388, 328, 516, 518, 520, 522, 404, 212, -1, -1, 524, 216, -1, -1, 526, 220, 528, 530, -1, -1, 532, 226, -1, -1, 534, 300, -1, -1, 536, 234, 538, 540, 456, 238, -1, -1, 542, 242, -1, -1, 544, 246, -1, -1, 546, 548, 550, 552, -1, -1, 554, 256, -1, -1, -1, -1, 262, 556, -1, -1, -1, -1, 558, 268, 270, 348, 560, 272, 274, 562, -1, -1, -1, -1, -1, -1, 282, 360, -1, -1, 564, 286, 288, 566, -1, -1, -1, -1, 294, 568, -1, -1, 298, 570, -1, -1, -1, -1, 412, 304, -1, -1, 308, 458, 354, 310, 312, 572, 314, 574, 576, 578, 580, 582, 584, 586, 588, 590, 466, 324, 326, 592, 368, 594, -1, -1, -1, -1, 596, 334, 598, 336, -1, -1, -1, -1, 342, 470, 346, 344, -1, -1, -1, -1, 350, 600, 602, 352, -1, -1, 604, 356, 606, 608, 610, 364, -1, -1, -1, -1, 366, 612, -1, -1, -1, -1, -1, -1, 614, 374, -1, -1, -1, -1, 380, 616, 384, 382, -1, -1, -1, -1, 618, 620, -1, -1, 622, 624, -1, -1, 626, 396, 628, 630, -1, -1, 452, 402, 632, 634, -1, -1, 474, 408, 410, 636, 482, 638, -1, -1, 416, 640, 642, 644, 646, 420, -1, -1, 648, 424, 650, 652, 654, 428, 656, 430, -1, -1, 658, 434, -1, -1, -1, -1, 440, 660, 662, 664, 478, 444, 666, 668, -1, -1, 670, 450, 672, 674, 454, 676, -1, -1, -1, -1, 460, 678, 680, 462, 464, 682, 684, 686, 468, 688, 690, 692, 472, 694, -1, -1, 696, 476, 698, 700, 702, 480, 704, 706, 708, 710, -1, -1, 712, 714, 716, 718, 720, 722, -1, -1, -1, -1, 724, 726, -1, -1, -1, -1, 728, 730, -1, -1, 732, 734, -1, -1, 736, 738, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 740, 742, -1, -1, -1, -1, -1, -1, -1, -1, 744, 746, 748, 750, 752, 754, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 756, 758, 760, 762, -1, -1, 764, 766, -1, -1, -1, -1, -1, -1, 768, 770, 772, 774, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 776, 778, -1, -1, 780, 782, -1, -1, 784, 786, -1, -1, 788, 790, 792, 794, 796, 798, 800, 802, -1, -1, -1, -1, 804, 806, -1, -1, -1, -1, -1, -1, -1, -1, 808, 810, -1, -1, -1, -1, -1, -1, -1, -1, 812, 814, 816, 818, 820, 822, -1, -1, -1, -1, -1, -1, 824, 826, -1, -1, -1, -1, 828, 830, -1, -1, -1, -1, 832, 834, -1, -1, -1, -1, 836, 838, 840, 842, 844, 846, -1, -1, -1, -1, -1, -1, 848, 850, 852, 854, 856, 858, -1, -1, -1, -1, 860, 862, -1, -1, -1, -1, -1, -1, 864, 866, 868, 870, 872, 874, 876, 878, -1, -1, -1, -1, -1, -1, -1, -1, 880, 882, 884, 886, 888, 890, 892, 894, 896, 898, 900, 902, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 952, 954, 956, 958, 960, 962, 964, 966, -1, -1, -1, -1, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, 14, 16, 18, 20, 12, 22, 24, 26, 28, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90, 92, 94, 96, 98, 100, 102, 104, 106, 108, 110, 112, 114, 116, 118, 120, 122, 124, 126, 128, 130, 132, 134, 136, 138, 140, 142, 144, 146, 148, 150, 152, 154, 156, 158, 160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 180, 182, 184, 186, 188, 190, 192, 194, 196, 198, 200, 202, 204, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, 432, 434, 436, 438, 440, 442, 444, 446, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, 512, 514, 516, 518, 520, 522, 524, 526, 528, 530, 532, 534, 536, 538, 540, 542, 544, 546, 548, 550, 552, 554, 556, 558, 560, 562, 564, 566, 568, 570, 572, 574, 576, 578, 580, 582, 584, 586, 588, 590, 592, 594, 596, 598, 600, 602, 604, 606, 608, 610, 612, 614, 616, 618, 620, 622, 624, 626, 628, 630, 632, 634, 636, 638, 640, 642, 644, 646, 648, 650, 652, 654, 656, 658, 660, 662, 664, 666, 668, 670, 672, 674, 676, 678, 680, 682, 684, 686, 688, 690, 692, 694, 696, 698, 700, 702, 704, 706, 708, 710, 712, 714, 716, 718, 720, 722, 724, 726, 728, 730, 732, 734, 736, 738, 740, 742, 744, 746, 748, 750, 752, 754, 756, 758, 760, 762, 764, 766, 768, 770, 772, 774, 776, 778, 780, 782, 784, 786, 788, 790, 792, 794, 796, 798, 800, 802, 804, 806, 808, 810, 812, 814, 816, 818, 820, 822, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 850, 852, 854, 856, 858, 860, 862, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, 888, 890, 892, 894, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 896, 898, 900, 902, 904, 906, 908, 910, 912, 914, 916, 918, 920, 922, 924, 926, 928, 930, 932, 934, 936, 938, 940, 942, 944, 946, 948, 950, 952, 954, 956, 958, 960, 962, 964, 966, 968, 970, 972, 974, 976, 978, 980, 982, 984, 986, 988, 990, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 10, 10, 5, 5, 4, 4, 16, 16, 13, 13, 12, 12, 6, 6, 24, 24, 11, 11, 27, 27, 21, 21, 30, 30, 17, 17, 35, 35, 9, 9, 40, 40, 41, 41, 22, 22, 46, 46, 8, 8, 49, 49, 52, 52, 15, 15, 55, 55, 58, 58, 14, 14, 61, 61, 19, 19, 65, 65, 18, 18, 69, 69, 53, 53, 74, 74, 47, 47, 72, 72, 20, 20, 81, 81, 26, 26, 85, 85, 87, 87, 75, 75, 32, 32, 93, 93, 25, 25, 98, 98, 96, 96, 29, 29, 104, 104, 80, 80, 31, 31, 109, 109, 99, 99, 113, 113, 37, 37, 117, 117, 106, 106, 44, 44, 123, 123, 33, 33, 64, 64, 125, 125, 34, 34, 133, 133, 79, 79, 78, 78, 57, 57, 142, 142, 129, 129, 43, 43, 148, 148, 149, 149, 137, 137, 60, 60, 108, 108, 89, 89, 38, 38, 162, 162, 105, 105, 23, 23, 167, 167, 170, 170, 128, 128, 145, 145, 28, 28, 178, 178, 163, 163, 36, 36, 184, 184, 185, 185, 171, 171, 189, 189, 111, 111, 76, 76, 112, 112, 144, 144, 91, 91, 82, 82, 179, 179, 90, 90, 42, 42, 209, 209, 211, 211, 56, 56, 215, 215, 218, 218, 220, 220, 221, 221, 73, 73, 225, 225, 59, 59, 84, 84, 232, 232, 54, 54, 235, 235, 237, 237, 62, 62, 242, 242, 92, 92, 50, 50, 247, 247, 250, 250, 51, 51, 254, 254, 255, 255, 155, 155, 259, 259, 203, 203, 264, 264, 86, 86, 267, 267, 269, 269, 251, 251, 274, 274, 83, 83, 107, 107, 97, 97, 39, 39, 284, 284, 285, 285, 288, 288, 289, 289, 287, 287, 138, 138, 77, 77, 48, 48, 63, 63, 302, 302, 195, 195, 172, 172, 187, 187, 258, 258, 100, 100, 45, 45, 315, 315, 318, 318, 281, 281, 88, 88, 120, 120, 150, 150, 239, 239, 214, 214, 126, 126, 188, 188, 227, 227, 217, 217, 340, 340, 124, 124, 344, 344, 134, 134, 169, 169, 350, 350, 177, 177, 354, 354, 356, 356, 249, 249, 360, 360, 361, 361, 94, 94, 366, 366, 127, 127, 238, 238, 371, 371, 252, 252, 375, 375, 161, 161, 380, 380, 180, 180, 383, 383, 230, 230, 387, 387, 226, 226, 391, 391, 299, 299, 241, 241, 398, 398, 210, 210, 402, 402, 216, 216, 405, 405, 408, 408, 406, 406, 412, 412, 70, 70, 415, 415, 283, 283, 420, 420, 66, 66, 67, 67, 68, 68, 71, 71, 95, 95, 103, 103, 110, 110, 114, 114, 118, 118, 119, 119, 130, 130, 141, 141, 143, 143, 146, 146, 147, 147, 156, 156, 164, 164, 168, 168, 183, 183, 186, 186, 190, 190, 196, 196, 199, 199, 200, 200, 204, 204, 205, 205, 206, 206, 212, 212, 213, 213, 219, 219, 222, 222, 228, 228, 229, 229, 231, 231, 236, 236, 240, 240, 243, 243, 244, 244, 248, 248, 253, 253, 256, 256, 257, 257, 260, 260, 263, 263, 268, 268, 270, 270, 273, 273, 275, 275, 276, 276, 277, 277, 278, 278, 282, 282, 286, 286, 290, 290, 293, 293, 294, 294, 300, 300, 301, 301, 303, 303, 304, 304, 307, 307, 308, 308, 311, 311, 312, 312, 313, 313, 314, 314, 316, 316, 317, 317, 321, 321, 322, 322, 323, 323, 324, 324, 339, 339, 341, 341, 342, 342, 343, 343, 349, 349, 351, 351, 352, 352, 353, 353, 355, 355, 359, 359, 362, 362, 363, 363, 364, 364, 365, 365, 372, 372, 376, 376, 377, 377, 378, 378, 379, 379, 384, 384, 388, 388, 392, 392, 397, 397, 399, 399, 400, 400, 401, 401, 403, 403, 404, 404, 407, 407, 409, 409, 410, 410, 411, 411, 413, 413, 414, 414, 416, 416, 417, 417, 418, 418, 419, 419, 421, 421, 422, 422, 423, 423, 424, 424, 425, 425, 426, 426, 427, 427, 428, 428, 429, 429, 430, 430, 433, 433, 434, 434, 435, 435, 436, 436, 439, 439, 440, 440, 443, 443, 444, 444, 445, 445, 446, 446, 447, 447, 448, 448, 451, 451, 452, 452, 453, 453, 454, 454, 457, 457, 458, 458, 459, 459, 460, 460, 461, 461, 462, 462, 471, 471, 472, 472, 477, 477, 478, 478, 481, 481, 482, 482, 487, 487, 488, 488, 491, 491, 492, 492, 495, 495, 496, 496, 497, 497, 498, 498, 499, 499, 500, 500, 501, 501, 502, 502, 503, 503, 504, 504, 505, 505, 506, 506, 511, 511, 512, 512, 515, 515, 516, 516, 525, 525, 526, 526, 527, 527, 528, 528, 537, 537, 538, 538, 555, 555, 556, 556, 567, 567, 568, 568, 575, 575, 576, 576, 581, 581, 582, 582, 585, 585, 586, 586, 587, 587, 588, 588, 597, 597, 598, 598, 611, 611, 612, 612, 617, 617, 618, 618, 623, 623, 624, 624, 629, 629, 630, 630, 635, 635, 636, 636, 637, 637, 638, 638, 639, 639, 640, 640, 641, 641, 642, 642, 643, 643, 644, 644, 645, 645, 646, 646, 647, 647, 648, 648, 649, 649, 650, 650, 659, 659, 660, 660, 661, 661, 662, 662, 679, 679, 680, 680, 681, 681, 682, 682, 695, 695, 696, 696, 697, 697, 698, 698, 699, 699, 700, 700, 701, 701, 702, 702, 723, 723, 724, 724, 725, 725, 726, 726, 735, 735, 736, 736, 737, 737, 738, 738, 739, 739, 740, 740, 741, 741, 742, 742, 743, 743, 744, 744, 745, 745, 746, 746, 763, 763, 764, 764, 765, 765, 766, 766, 787, 787, 788, 788, 789, 789, 790, 790, 815, 815, 816, 816, 817, 817, 818, 818, 827, 827, 828, 828, 829, 829, 830, 830, 863, 863, 864, 864, 865, 865, 866, 866, 867, 867, 868, 868, 869, 869, 870, 870, 887, 887, 888, 888, 889, 889, 890, 890, 891, 891, 892, 892, 893, 893, 894, 894, 895, 895, 896, 896, 897, 897, 898, 898, 899, 899, 900, 900, 901, 901, 902, 902, 959, 959, 960, 960, 961, 961, 962, 962, 963, 963, 964, 964, 965, 965, 966, 966, 967, 967, 968, 968, 969, 969, 970, 970, 971, 971, 972, 972, 973, 973, 974, 974),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 10, 10, 4, 4, 14, 14, 5, 5, 17, 17, 6, 6, 21, 21, 16, 16, 26, 26, 15, 15, 27, 27, 30, 30, 11, 11, 35, 35, 12, 12, 39, 39, 9, 9, 44, 44, 33, 33, 45, 45, 18, 18, 52, 52, 37, 37, 42, 42, 8, 8, 59, 59, 62, 62, 48, 48, 13, 13, 67, 67, 70, 70, 38, 38, 31, 31, 19, 19, 77, 77, 63, 63, 56, 56, 82, 82, 24, 24, 71, 71, 90, 90, 83, 83, 65, 65, 36, 36, 98, 98, 100, 100, 28, 28, 104, 104, 51, 51, 107, 107, 25, 25, 111, 111, 114, 114, 58, 58, 32, 32, 120, 120, 46, 46, 123, 123, 29, 29, 128, 128, 129, 129, 130, 130, 61, 61, 136, 136, 20, 20, 139, 139, 73, 73, 84, 84, 137, 137, 23, 23, 150, 150, 125, 125, 102, 102, 88, 88, 69, 69, 160, 160, 53, 53, 164, 164, 89, 89, 168, 168, 22, 22, 171, 171, 174, 174, 54, 54, 177, 177, 75, 75, 118, 118, 148, 148, 133, 133, 49, 49, 190, 190, 92, 92, 57, 57, 195, 195, 76, 76, 87, 87, 202, 202, 142, 142, 152, 152, 86, 86, 210, 210, 161, 161, 214, 214, 173, 173, 218, 218, 153, 153, 80, 80, 224, 224, 110, 110, 106, 106, 40, 40, 232, 232, 103, 103, 236, 236, 99, 99, 240, 240, 47, 47, 244, 244, 79, 79, 158, 158, 192, 192, 162, 162, 254, 254, 131, 131, 74, 74, 259, 259, 180, 180, 68, 68, 266, 266, 267, 267, 270, 270, 271, 271, 116, 116, 143, 143, 85, 85, 279, 279, 72, 72, 284, 284, 285, 285, 66, 66, 55, 55, 291, 291, 175, 175, 295, 295, 228, 228, 113, 113, 302, 302, 60, 60, 305, 305, 308, 308, 309, 309, 311, 311, 126, 126, 141, 141, 163, 163, 172, 172, 322, 322, 323, 323, 204, 204, 91, 91, 149, 149, 332, 332, 334, 334, 154, 154, 112, 112, 339, 339, 342, 342, 341, 341, 268, 268, 347, 347, 350, 350, 307, 307, 354, 354, 81, 81, 280, 280, 167, 167, 358, 358, 363, 363, 325, 325, 165, 165, 109, 109, 372, 372, 144, 144, 97, 97, 377, 377, 380, 380, 379, 379, 157, 157, 203, 203, 147, 147, 105, 105, 78, 78, 394, 394, 101, 101, 108, 108, 400, 400, 209, 209, 43, 43, 406, 406, 407, 407, 301, 301, 138, 138, 413, 413, 201, 201, 418, 418, 41, 41, 422, 422, 159, 159, 426, 426, 428, 428, 178, 178, 432, 432, 179, 179, 124, 124, 437, 437, 135, 135, 442, 442, 119, 119, 140, 140, 448, 448, 399, 399, 451, 451, 235, 235, 306, 306, 457, 457, 460, 460, 461, 461, 321, 321, 465, 465, 340, 340, 469, 469, 405, 405, 474, 474, 441, 441, 478, 478, 409, 409, 186, 186, 34, 34, 50, 50, 64, 64, 115, 115, 117, 117, 127, 127, 132, 132, 134, 134, 151, 151, 166, 166, 176, 176, 185, 185, 189, 189, 191, 191, 196, 196, 205, 205, 206, 206, 207, 207, 208, 208, 213, 213, 217, 217, 219, 219, 220, 220, 223, 223, 227, 227, 231, 231, 233, 233, 234, 234, 239, 239, 243, 243, 247, 247, 248, 248, 249, 249, 250, 250, 253, 253, 260, 260, 265, 265, 269, 269, 272, 272, 283, 283, 286, 286, 292, 292, 296, 296, 310, 310, 312, 312, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 318, 318, 319, 319, 320, 320, 324, 324, 326, 326, 331, 331, 333, 333, 348, 348, 349, 349, 353, 353, 355, 355, 356, 356, 357, 357, 364, 364, 371, 371, 378, 378, 385, 385, 386, 386, 389, 389, 390, 390, 393, 393, 395, 395, 396, 396, 401, 401, 402, 402, 408, 408, 410, 410, 414, 414, 415, 415, 416, 416, 417, 417, 421, 421, 423, 423, 424, 424, 425, 425, 427, 427, 431, 431, 438, 438, 439, 439, 440, 440, 443, 443, 444, 444, 447, 447, 449, 449, 450, 450, 452, 452, 458, 458, 459, 459, 462, 462, 463, 463, 464, 464, 466, 466, 467, 467, 468, 468, 470, 470, 473, 473, 475, 475, 476, 476, 477, 477, 479, 479, 480, 480, 481, 481, 482, 482, 485, 485, 486, 486, 487, 487, 488, 488, 489, 489, 490, 490, 495, 495, 496, 496, 501, 501, 502, 502, 505, 505, 506, 506, 509, 509, 510, 510, 525, 525, 526, 526, 535, 535, 536, 536, 537, 537, 538, 538, 539, 539, 540, 540, 557, 557, 558, 558, 559, 559, 560, 560, 563, 563, 564, 564, 571, 571, 572, 572, 573, 573, 574, 574, 591, 591, 592, 592, 595, 595, 596, 596, 599, 599, 600, 600, 603, 603, 604, 604, 605, 605, 606, 606, 607, 607, 608, 608, 609, 609, 610, 610, 615, 615, 616, 616, 625, 625, 626, 626, 635, 635, 636, 636, 637, 637, 638, 638, 639, 639, 640, 640, 647, 647, 648, 648, 653, 653, 654, 654, 659, 659, 660, 660, 665, 665, 666, 666, 667, 667, 668, 668, 669, 669, 670, 670, 677, 677, 678, 678, 679, 679, 680, 680, 681, 681, 682, 682, 687, 687, 688, 688, 695, 695, 696, 696, 697, 697, 698, 698, 699, 699, 700, 700, 701, 701, 702, 702, 711, 711, 712, 712, 713, 713, 714, 714, 715, 715, 716, 716, 717, 717, 718, 718, 719, 719, 720, 720, 721, 721, 722, 722, 723, 723, 724, 724, 725, 725, 726, 726, 743, 743, 744, 744, 745, 745, 746, 746, 755, 755, 756, 756, 757, 757, 758, 758, 767, 767, 768, 768, 769, 769, 770, 770, 787, 787, 788, 788, 789, 789, 790, 790, 811, 811, 812, 812, 813, 813, 814, 814, 847, 847, 848, 848, 849, 849, 850, 850, 851, 851, 852, 852, 853, 853, 854, 854, 863, 863, 864, 864, 865, 865, 866, 866, 895, 895, 896, 896, 897, 897, 898, 898, 899, 899, 900, 900, 901, 901, 902, 902, 919, 919, 920, 920, 921, 921, 922, 922, 923, 923, 924, 924, 925, 925, 926, 926, 951, 951, 952, 952, 953, 953, 954, 954, 955, 955, 956, 956, 957, 957, 958, 958),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 10, 10, 11, 11, 12, 12, 13, 13, 14, 14, 15, 15, 16, 16, 17, 17, 18, 18, 19, 19, 20, 20, 21, 21, 22, 22, 23, 23, 24, 24, 25, 25, 26, 26, 27, 27, 28, 28, 29, 29, 30, 30, 31, 31, 32, 32, 33, 33, 34, 34, 35, 35, 36, 36, 37, 37, 38, 38, 39, 39, 40, 40, 41, 41, 42, 42, 43, 43, 44, 44, 45, 45, 46, 46, 47, 47, 48, 48, 49, 49, 50, 50, 51, 51, 52, 52, 53, 53, 54, 54, 55, 55, 56, 56, 57, 57, 58, 58, 59, 59, 60, 60, 61, 61, 62, 62, 63, 63, 64, 64, 65, 65, 66, 66, 67, 67, 68, 68, 69, 69, 70, 70, 71, 71, 72, 72, 73, 73, 74, 74, 75, 75, 76, 76, 77, 77, 78, 78, 79, 79, 80, 80, 81, 81, 82, 82, 83, 83, 84, 84, 85, 85, 86, 86, 87, 87, 88, 88, 89, 89, 90, 90, 91, 91, 92, 92, 93, 93, 94, 94, 95, 95, 96, 96, 97, 97, 98, 98, 99, 99, 100, 100, 101, 101, 102, 102, 103, 103, 104, 104, 105, 105, 106, 106, 107, 107, 108, 108, 109, 109, 110, 110, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 117, 117, 118, 118, 119, 119, 120, 120, 121, 121, 122, 122, 123, 123, 124, 124, 125, 125, 126, 126, 127, 127, 128, 128, 129, 129, 130, 130, 131, 131, 132, 132, 133, 133, 134, 134, 135, 135, 136, 136, 137, 137, 138, 138, 139, 139, 140, 140, 141, 141, 142, 142, 143, 143, 144, 144, 145, 145, 146, 146, 147, 147, 148, 148, 149, 149, 150, 150, 151, 151, 152, 152, 153, 153, 154, 154, 155, 155, 156, 156, 157, 157, 158, 158, 159, 159, 160, 160, 161, 161, 162, 162, 163, 163, 164, 164, 165, 165, 166, 166, 167, 167, 168, 168, 169, 169, 170, 170, 171, 171, 172, 172, 173, 173, 174, 174, 175, 175, 176, 176, 177, 177, 178, 178, 179, 179, 180, 180, 181, 181, 182, 182, 183, 183, 184, 184, 185, 185, 186, 186, 187, 187, 188, 188, 189, 189, 190, 190, 191, 191, 192, 192, 193, 193, 194, 194, 195, 195, 196, 196, 197, 197, 198, 198, 199, 199, 200, 200, 201, 201, 202, 202, 203, 203, 204, 204, 205, 205, 206, 206, 207, 207, 208, 208, 209, 209, 210, 210, 211, 211, 212, 212, 213, 213, 214, 214, 215, 215, 216, 216, 217, 217, 218, 218, 219, 219, 220, 220, 221, 221, 222, 222, 223, 223, 224, 224, 225, 225, 226, 226, 227, 227, 228, 228, 229, 229, 230, 230, 231, 231, 232, 232, 233, 233, 234, 234, 235, 235, 236, 236, 237, 237, 238, 238, 239, 239, 240, 240, 241, 241, 242, 242, 243, 243, 244, 244, 245, 245, 246, 246, 247, 247, 248, 248, 249, 249, 250, 250, 251, 251, 252, 252, 253, 253, 254, 254, 255, 255, 256, 256, 257, 257, 258, 258, 259, 259, 260, 260, 261, 261, 262, 262, 263, 263, 264, 264, 265, 265, 266, 266, 267, 267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 272, 273, 273, 274, 274, 275, 275, 276, 276, 277, 277, 278, 278, 279, 279, 280, 280, 281, 281, 282, 282, 283, 283, 284, 284, 285, 285, 286, 286, 287, 287, 288, 288, 289, 289, 290, 290, 291, 291, 292, 292, 293, 293, 294, 294, 295, 295, 296, 296, 297, 297, 298, 298, 299, 299, 300, 300, 301, 301, 302, 302, 303, 303, 304, 304, 305, 305, 306, 306, 307, 307, 308, 308, 309, 309, 310, 310, 311, 311, 312, 312, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 323, 323, 324, 324, 325, 325, 326, 326, 327, 327, 328, 328, 329, 329, 330, 330, 331, 331, 332, 332, 333, 333, 334, 334, 335, 335, 336, 336, 337, 337, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 345, 345, 346, 346, 347, 347, 348, 348, 349, 349, 350, 350, 351, 351, 352, 352, 353, 353, 354, 354, 355, 355, 356, 356, 357, 357, 358, 358, 359, 359, 360, 360, 361, 361, 362, 362, 363, 363, 364, 364, 365, 365, 366, 366, 367, 367, 368, 368, 369, 369, 370, 370, 371, 371, 372, 372, 373, 373, 374, 374, 375, 375, 376, 376, 377, 377, 378, 378, 379, 379, 380, 380, 381, 381, 382, 382, 383, 383, 384, 384, 385, 385, 386, 386, 387, 387, 388, 388, 389, 389, 390, 390, 391, 391, 392, 392, 393, 393, 394, 394, 395, 395, 396, 396, 397, 397, 398, 398, 399, 399, 400, 400, 401, 401, 402, 402, 403, 403, 404, 404, 405, 405, 406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 412, 412, 413, 413, 414, 414, 415, 415, 416, 416, 417, 417, 418, 418, 419, 419, 420, 420, 421, 421, 422, 422, 423, 423, 424, 424, 425, 425, 426, 426, 427, 427, 428, 428, 429, 429, 430, 430, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446, 703, 703, 704, 704, 705, 705, 706, 706, 707, 707, 708, 708, 709, 709, 710, 710, 711, 711, 712, 712, 713, 713, 714, 714, 715, 715, 716, 716, 717, 717, 718, 718, 719, 719, 720, 720, 721, 721, 722, 722, 723, 723, 724, 724, 725, 725, 726, 726, 727, 727, 728, 728, 729, 729, 730, 730, 731, 731, 732, 732, 733, 733, 734, 734, 735, 735, 736, 736, 737, 737, 738, 738, 739, 739, 740, 740, 741, 741, 742, 742, 743, 743, 744, 744, 745, 745, 746, 746, 747, 747, 748, 748, 749, 749, 750, 750, 751, 751, 752, 752, 753, 753, 754, 754, 755, 755, 756, 756, 757, 757, 758, 758, 759, 759, 760, 760, 761, 761, 762, 762, 763, 763, 764, 764, 765, 765, 766, 766)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 3, 3, 4, 4, 5, 5, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 7, 7, 5, 5, 6, 6, 4, 4, 5, 5, 6, 6, 6, 6, 7, 7, 3, 3, 4, 4, 5, 5, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 6, 6, 7, 7, 5, 5, 6, 6, 6, 6, 7, 7, 8, 8, 7, 7, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 9, 9, 9, 9, 6, 6, 7, 7, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 9, 9, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 9, 9, 8, 8, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 3, 3, 4, 4, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 5, 5, 7, 7, 6, 6, 5, 5, 6, 6, 5, 5, 6, 6, 4, 4, 5, 5, 7, 7, 6, 6, 5, 5, 6, 6, 7, 7, 7, 7, 3, 3, 4, 4, 5, 5, 8, 8, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 8, 8, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 5, 5, 6, 6, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 6, 6, 7, 7, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 7, 7, 6, 6, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 6, 6, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((101, 102, 115, 116, 121, 122, 131, 132, 135, 136, 139, 140, 151, 152, 153, 154, 157, 158, 159, 160, 165, 166, 173, 174, 175, 176, 181, 182, 191, 192, 193, 194, 197, 198, 201, 202, 207, 208, 223, 224, 233, 234, 245, 246, 261, 262, 265, 266, 271, 272, 279, 280, 291, 292, 295, 296, 297, 298, 305, 306, 309, 310, 319, 320, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 345, 346, 347, 348, 357, 358, 367, 368, 369, 370, 373, 374, 381, 382, 385, 386, 389, 390, 393, 394, 395, 396, 431, 432, 437, 438, 441, 442, 449, 450, 455, 456, 463, 464, 465, 466, 467, 468, 469, 470, 473, 474, 475, 476, 479, 480, 483, 484, 485, 486, 489, 490, 493, 494, 507, 508, 509, 510, 513, 514, 517, 518, 519, 520, 521, 522, 523, 524, 529, 530, 531, 532, 533, 534, 535, 536, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 569, 570, 571, 572, 573, 574, 577, 578, 579, 580, 583, 584, 589, 590, 591, 592, 593, 594, 595, 596, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 613, 614, 615, 616, 619, 620, 621, 622, 625, 626, 627, 628, 631, 632, 633, 634, 651, 652, 653, 654, 655, 656, 657, 658, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 727, 728, 729, 730, 731, 732, 733, 734, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 759, 760, 761, 762, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 819, 820, 821, 822, 823, 824, 825, 826, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (93, 94, 95, 96, 121, 122, 145, 146, 155, 156, 169, 170, 181, 182, 183, 184, 187, 188, 193, 194, 197, 198, 199, 200, 211, 212, 215, 216, 221, 222, 225, 226, 229, 230, 237, 238, 241, 242, 245, 246, 251, 252, 255, 256, 257, 258, 261, 262, 263, 264, 273, 274, 275, 276, 277, 278, 281, 282, 287, 288, 289, 290, 293, 294, 297, 298, 299, 300, 303, 304, 327, 328, 329, 330, 335, 336, 337, 338, 343, 344, 345, 346, 351, 352, 359, 360, 361, 362, 365, 366, 367, 368, 369, 370, 373, 374, 375, 376, 381, 382, 383, 384, 387, 388, 391, 392, 397, 398, 403, 404, 411, 412, 419, 420, 429, 430, 433, 434, 435, 436, 445, 446, 453, 454, 455, 456, 471, 472, 483, 484, 491, 492, 493, 494, 497, 498, 499, 500, 503, 504, 507, 508, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 527, 528, 529, 530, 531, 532, 533, 534, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 561, 562, 565, 566, 567, 568, 569, 570, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 593, 594, 597, 598, 601, 602, 611, 612, 613, 614, 617, 618, 619, 620, 621, 622, 623, 624, 627, 628, 629, 630, 631, 632, 633, 634, 641, 642, 643, 644, 645, 646, 649, 650, 651, 652, 655, 656, 657, 658, 661, 662, 663, 664, 671, 672, 673, 674, 675, 676, 683, 684, 685, 686, 689, 690, 691, 692, 693, 694, 703, 704, 705, 706, 707, 708, 709, 710, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 747, 748, 749, 750, 751, 752, 753, 754, 759, 760, 761, 762, 763, 764, 765, 766, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 855, 856, 857, 858, 859, 860, 861, 862, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 863, 864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
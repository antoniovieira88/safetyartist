library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((2, 2, 1, 1, 1, 1, 0, -2, -2, 1, -2, -2, 1, -2, 1, -2, -2, 0, 0, -2, 0, -2, -2, 1, 1, -2, -2, 0, -2, -2, 1, 0, 1, 0, -2, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 0, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 0, 2, 0, 0, 0, -2, -2, 1, -2, -2, 0, 1, -2, -2, 0, -2, -2, 1, 1, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, 1, -2, -2, 2, 0, 1, 0, -2, -2, 1, -2, -2, 1, 1, -2, -2, 0, -2, -2, 1, 0, 1, -2, -2, 1, -2, -2, 0, 1, -2, -2, 1, -2, -2, 2, 1, 0, 1, 1, 0, -2, -2, 0, -2, -2, 1, 1, -2, -2, -2, 0, 1, 1, -2, -2, 1, -2, -2, 0, 1, -2, -2, -2, 1, 1, -2, 0, 1, -2, -2, 0, -2, -2, 1, 0, 1, -2, -2, 1, -2, -2, -2, 0, 1, 0, 1, 0, -2, -2, 0, -2, -2, 1, 1, -2, -2, 0, -2, -2, 1, 0, -2, 0, -2, -2, 1, 0, -2, -2, -2, 0, 1, 0, 1, -2, -2, 1, -2, -2, 1, 0, -2, -2, -2, 1, -2, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 2, 0, 0, 0, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 0, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, -2, 1, 0, 0, -2, 0, -2, -2, 1, 2, -2, -2, 0, -2, -2, 2, 0, 0, -2, -2, 1, -2, -2, 0, 1, -2, -2, 0, -2, -2, 1, 1, 2, 1, 0, -2, -2, 0, -2, -2, 1, -2, 2, -2, -2, 1, 1, -2, 1, -2, -2, 2, 1, -2, -2, 2, -2, -2, 1, 2, 1, 1, -2, -2, 1, -2, -2, 1, -2, 1, -2, -2, 1, -2, 2, 1, -2, -2, 0, -2, -2, 0, 1, 1, 1, 0, -2, -2, 0, 2, -2, -2, 1, -2, -2, 1, 0, -2, -2, 2, 1, -2, -2, 0, -2, -2, 2, 0, 0, 0, -2, -2, 1, -2, -2, 1, 1, -2, -2, -2, 0, 1, 0, -2, -2, 1, -2, -2, 1, 1, -2, -2, 1, -2, -2, 2, 0, 0, 0, 1, -2, -2, 1, -2, -2, 1, 1, -2, -2, 0, -2, -2, 0, 1, 0, -2, -2, 1, -2, -2, -2, 0, 0, 0, -2, 0, -2, -2, -2, 0, 1, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 2, 1, 1, 1, 0, -2, -2, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, 1, 0, 1, -2, -2, 0, -2, -2, 1, 1, -2, -2, -2, 1, 1, 0, 2, -2, -2, 2, -2, -2, 0, 2, -2, -2, 2, -2, -2, 1, 1, 0, -2, -2, 1, -2, -2, 2, 1, -2, -2, 0, -2, -2, 0, 2, 0, 1, 0, -2, -2, 0, -2, -2, 1, 1, -2, -2, 1, -2, -2, 1, 1, 0, -2, -2, 0, -2, -2, 1, 0, -2, -2, -2, 0, 1, 1, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, 2, -2, -2, 1, 2, 0, -2, -2, 0, -2, -2, 1, 2, -2, -2, 1, -2, -2, 1, 1, 1, 0, 1, -2, 2, -2, -2, -2, 0, 0, 2, -2, -2, 2, -2, -2, 2, 0, -2, -2, 2, -2, -2, 0, 2, 2, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 2, 0, 1, -2, -2, -2, 0, 1, -2, -2, -2, 1, 2, 0, 0, 1, -2, -2, 1, -2, -2, 0, 0, -2, -2, -2, 1, -2, 0, 0, -2, -2, 0, -2, -2, 0, 1, 1, 2, -2, -2, -2, 2, 1, -2, -2, 0, -2, -2, 1, 1, -2, 0, -2, -2, 0, 2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((134, 92, 2228, 1736, 768, 593, 1980, -256, -256, 594, -256, -256, 770, -256, 899, -256, -256, 28048, 26709, -256, 27089, -256, -256, 2044, 1979, -256, -256, 35806, -256, -256, 2948, 49942, 2418, 41192, -256, -256, -256, 56522, 2790, -256, -256, 2805, -256, -256, 74130, 66599, 2997, -256, -256, 66600, -256, -256, 80935, 3233, -256, -256, 88178, -256, -256, 38395, 109, 19001, 5007, 3874, -256, -256, 1305, -256, -256, 30769, 1803, -256, -256, 38054, -256, -256, 1835, 889, 765, -256, -256, 1497, -256, -256, 33138, 25321, -256, -256, 2651, -256, -256, 109, 63871, 2918, 47283, -256, -256, 3085, -256, -256, 3461, 3330, -256, -256, 74797, -256, -256, 2886, 38480, 2196, -256, -256, 2790, -256, -256, 60065, 3313, -256, -256, 3461, -256, -256, 164, 2187, 12856, 971, 384, 632, -256, -256, 3736, -256, -256, 1341, 1314, -256, -256, -256, 20604, 1815, 1649, -256, -256, 1902, -256, -256, 23014, 2067, -256, -256, -256, 2940, 2188, -256, 31705, 2237, -256, -256, 34761, -256, -256, 3798, 48932, 3063, -256, -256, 3460, -256, -256, -256, 23282, 1549, 3685, 329, 612, -256, -256, 2738, -256, -256, 1087, 856, -256, -256, 11672, -256, -256, 1992, 15398, -256, 16572, -256, -256, 2181, 20650, -256, -256, -256, 38339, 2541, 24138, 2140, -256, -256, 2472, -256, -256, 3107, 33107, -256, -256, -256, 3228, -256, 3228, -256, 3658, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256),
                (134, 2102, 92, 20559, 7992, 1305, 64, -256, -256, 1321, -256, -256, 15103, 1024, -256, -256, 1402, -256, -256, 28029, 27884, 1772, -256, -256, 27891, -256, -256, 33546, 2024, -256, -256, -256, 1264, 4796, 1150, -256, 3700, -256, -256, 930, 109, -256, -256, 10130, -256, -256, 109, 21732, 16443, -256, -256, 2010, -256, -256, 19366, 1563, -256, -256, 24495, -256, -256, 2808, 2404, 92, 2111, 32660, -256, -256, 37208, -256, -256, 2102, -256, 109, -256, -256, 2406, 2405, -256, 2405, -256, -256, 92, 2779, -256, -256, 109, -256, -256, 3033, 109, 3025, 3022, -256, -256, 3031, -256, -256, 2808, -256, 3026, -256, -256, 3033, -256, 92, 3288, -256, -256, 63950, -256, -256, 26703, 1453, 855, 193, 587, -256, -256, 2550, 164, -256, -256, 834, -256, -256, 876, 8208, -256, -256, 164, 1403, -256, -256, 9079, -256, -256, 164, 19098, 16490, 15208, -256, -256, 1803, -256, -256, 2240, 1933, -256, -256, -256, 16626, 1776, 12850, -256, -256, 1864, -256, -256, 2200, 2024, -256, -256, 2323, -256, -256, 164, 43118, 34496, 27968, 2248, -256, -256, 2602, -256, -256, 2878, 2744, -256, -256, 41980, -256, -256, 55317, 3224, 44806, -256, -256, 3467, -256, -256, -256, 35807, 35794, 26901, -256, 26993, -256, -256, -256, 46325, 3294, 37238, -256, -256, 41600, -256, -256, 47566, 3538, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256),
                (39757, 134, 92, 1728, 1190, 830, 3768, -256, -256, 1165, -256, -256, 1629, 15952, -256, -256, 1700, -256, -256, 2073, 27984, 1792, -256, -256, 31496, -256, -256, 2195, 2187, -256, -256, -256, 1677, 928, 3899, 109, -256, -256, 109, -256, -256, 13769, 109, -256, -256, 109, -256, -256, 2245, 1912, 20553, -256, -256, 2243, -256, -256, 109, 2578, -256, -256, 39588, -256, -256, 12852, 164, 3722, 254, 622, -256, -256, 2497, -256, -256, 1083, 881, -256, -256, 1342, -256, -256, 1067, 329, 1142, -256, -256, 3782, -256, -256, 1399, 9065, -256, -256, -256, 20576, 1768, 1632, 1416, -256, -256, 1665, -256, -256, 19477, 17261, -256, -256, 164, -256, -256, 2541, 164, 30563, -256, -256, 24138, -256, -256, 2941, 164, -256, -256, 3105, -256, -256, 2938, 2714, 2454, 44755, 2341, -256, 92, -256, -256, -256, 45761, 42059, 109, -256, -256, 92, -256, -256, 92, 49382, -256, -256, 109, -256, -256, 55090, 109, 92, 2754, -256, -256, 47368, -256, -256, 41886, 2801, -256, -256, 43541, -256, -256, 92, 62717, 2798, -256, -256, -256, 57541, 2918, -256, -256, -256, 3232, 109, 62703, 60424, 3016, -256, -256, 3119, -256, -256, 72788, 72747, -256, -256, -256, 2938, -256, 48298, 44670, -256, -256, 52175, -256, -256, 66440, 3403, 3402, 134, -256, -256, -256, 134, 3503, -256, -256, 48156, -256, -256, 3462, 3271, -256, 75724, -256, -256, 74110, 109, -256, -256, 92, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((38, 38, 37, 40, 41, 42, 42, 7, 43, 42, 0, 42, 40, 0, 40, 41, 40, 37, 1, 0, 9, 21, 0, 42, 43, 43, 42, 41, 3, 42, 32, 34, 2, 7, 0, 41, 0, 42, 28, 40, 0, 42, 43, 42, 30, 1, 0, 1, 0, 9, 43, 8, 42, 23, 43, 6, 42, 37, 43, 38, 18, 17, 10, 3, 2, 7, 13, 38, 1, 23, 21, 42, 2, 27, 28, 13, 18, 32, 39, 40, 34, 24, 27, 20, 4, 2, 0, 7, 20, 40, 0, 42, 42, 34, 41, 38, 42, 5, 17, 1, 43, 43, 43, 42, 40, 2, 43, 42, 43, 28, 43, 0, 43, 43, 42, 39, 7, 12, 1, 42, 43, 41, 39, 39, 41, 17, 34, 41, 0, 43, 27, 0, 38, 4, 14, 11, 30, 0, 42, 36, 42, 43, 30, 1, 4, 0, 43, 40, 43, 0, 43, 36, 38, 0, 38, 2, 14, 1, 42, 31, 43, 34, 34, 2, 7, 0, 42, 43, 41, 0, 39, 15, 31, 5, 18, 0, 38, 1, 0, 6, 38, 42, 43, 39, 28, 4, 43, 3, 14, 0, 41, 28, 43, 1, 5, 0, 43, 0, 42, 31, 42, 34, 43, 0, 42, 43, 35, 7, 14, 6, 30, 0, 43, 43, 41, 0, 41, 41, 39, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43),
                (38, 38, 41, 40, 19, 11, 1, 21, 0, 14, 43, 13, 26, 22, 42, 3, 30, 43, 3, 42, 36, 37, 42, 0, 9, 0, 21, 43, 41, 42, 5, 43, 41, 42, 10, 0, 14, 11, 22, 42, 43, 43, 43, 42, 5, 43, 39, 39, 4, 0, 16, 42, 43, 41, 39, 4, 11, 0, 42, 32, 43, 33, 36, 37, 35, 27, 0, 43, 36, 0, 42, 37, 0, 37, 37, 37, 35, 17, 0, 21, 43, 14, 35, 33, 33, 37, 35, 35, 36, 32, 33, 32, 32, 32, 18, 40, 42, 32, 34, 0, 34, 34, 43, 31, 0, 31, 29, 31, 28, 32, 2, 42, 39, 17, 34, 38, 41, 0, 43, 37, 2, 3, 0, 42, 42, 36, 28, 5, 0, 43, 29, 28, 27, 37, 29, 3, 42, 5, 5, 1, 0, 0, 1, 5, 43, 0, 15, 37, 43, 31, 0, 5, 1, 4, 0, 43, 0, 2, 0, 12, 37, 43, 27, 2, 13, 0, 42, 42, 32, 30, 35, 43, 0, 28, 41, 0, 34, 42, 43, 27, 1, 0, 11, 43, 41, 43, 42, 43, 16, 21, 0, 43, 42, 32, 32, 43, 32, 13, 32, 0, 43, 39, 42, 39, 42, 6, 0, 11, 43, 42, 43, 0, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0),
                (38, 20, 19, 17, 33, 37, 39, 9, 42, 33, 32, 43, 24, 25, 2, 41, 19, 16, 36, 2, 9, 1, 6, 0, 39, 32, 41, 0, 3, 2, 43, 0, 19, 34, 39, 15, 16, 15, 42, 42, 42, 28, 5, 5, 5, 41, 40, 42, 5, 15, 18, 0, 40, 13, 13, 43, 1, 1, 2, 0, 1, 1, 32, 22, 10, 10, 2, 38, 0, 43, 1, 0, 3, 13, 40, 41, 31, 2, 16, 0, 11, 31, 39, 7, 43, 28, 3, 41, 2, 10, 1, 43, 0, 28, 22, 42, 42, 43, 40, 30, 9, 36, 2, 1, 0, 2, 7, 5, 9, 31, 41, 40, 38, 43, 42, 38, 43, 5, 15, 8, 22, 1, 3, 0, 42, 43, 43, 43, 43, 43, 39, 0, 43, 43, 42, 31, 36, 19, 43, 27, 0, 41, 43, 42, 7, 43, 43, 43, 43, 41, 25, 7, 1, 6, 0, 13, 0, 24, 39, 24, 43, 20, 42, 39, 43, 42, 42, 24, 36, 17, 43, 43, 39, 43, 26, 43, 39, 40, 38, 3, 1, 4, 0, 21, 38, 0, 42, 32, 34, 0, 43, 42, 0, 42, 21, 16, 27, 42, 34, 43, 38, 13, 15, 15, 2, 35, 43, 11, 2, 3, 0, 27, 5, 39, 42, 42, 43, 42, 32, 43, 41, 24, 3, 43, 42, 40, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 3, 4, 5, 6, 7, -1, -1, 10, -1, -1, 13, 219, 15, -1, -1, 18, 19, 221, 21, -1, -1, 24, 25, -1, -1, 28, -1, -1, 31, 32, 33, 34, -1, -1, 223, 38, 39, -1, -1, 42, -1, -1, 45, 46, 47, -1, -1, 50, -1, -1, 53, 54, -1, -1, 57, -1, -1, 60, 61, 62, 63, 64, -1, -1, 67, -1, -1, 70, 71, -1, -1, 74, -1, -1, 77, 78, 79, -1, -1, 82, -1, -1, 85, 86, -1, -1, 89, -1, -1, 92, 93, 94, 95, -1, -1, 98, -1, -1, 101, 102, -1, -1, 105, -1, -1, 108, 109, 110, -1, -1, 113, -1, -1, 116, 117, -1, -1, 120, -1, -1, 123, 124, 125, 126, 127, 128, -1, -1, 131, -1, -1, 134, 135, -1, -1, 225, 139, 140, 141, -1, -1, 144, -1, -1, 147, 148, -1, -1, 227, 152, 153, 229, 155, 156, -1, -1, 159, -1, -1, 162, 163, 164, -1, -1, 167, -1, -1, 231, 171, 172, 173, 174, 175, -1, -1, 178, -1, -1, 181, 182, -1, -1, 185, -1, -1, 188, 189, 233, 191, -1, -1, 194, 195, -1, -1, 235, 199, 200, 201, 202, -1, -1, 205, -1, -1, 208, 209, -1, -1, 237, 213, 239, 215, 241, 217, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 243, 245, 247, 249, -1, -1, -1, -1, -1, -1, 251, 253, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, 7, -1, -1, 10, -1, -1, 13, 14, -1, -1, 17, -1, -1, 20, 21, 22, -1, -1, 25, -1, -1, 28, 29, -1, -1, 213, 33, 34, 35, 215, 37, -1, -1, 40, 41, -1, -1, 44, -1, -1, 47, 48, 49, -1, -1, 52, -1, -1, 55, 56, -1, -1, 59, -1, -1, 62, 63, 64, 65, 66, -1, -1, 69, -1, -1, 72, 217, 74, -1, -1, 77, 78, 219, 80, -1, -1, 83, 84, -1, -1, 87, -1, -1, 90, 91, 92, 93, -1, -1, 96, -1, -1, 99, 221, 101, -1, -1, 104, 223, 106, 107, -1, -1, 110, -1, -1, 113, 114, 115, 116, 117, 225, 227, 120, 121, -1, -1, 124, -1, -1, 127, 128, 229, 231, 131, 132, -1, -1, 135, -1, -1, 138, 139, 140, 141, -1, -1, 144, -1, -1, 147, 148, -1, -1, 233, 152, 153, 154, -1, -1, 157, -1, -1, 160, 161, -1, -1, 164, -1, -1, 167, 168, 169, 170, 171, -1, -1, 174, -1, -1, 177, 178, -1, -1, 181, -1, -1, 184, 185, 186, -1, -1, 189, -1, -1, 235, 193, 194, 195, 237, 197, -1, -1, 239, 201, 202, 203, -1, -1, 206, -1, -1, 209, 210, -1, -1, 241, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 243, 245, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 247, 249, -1, -1, 251, 253, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, 7, -1, -1, 10, -1, -1, 13, 14, -1, -1, 17, -1, -1, 20, 21, 22, -1, -1, 25, -1, -1, 28, 29, -1, -1, 227, 33, 34, 35, 36, -1, -1, 39, -1, -1, 42, 43, -1, -1, 46, -1, -1, 49, 50, 51, -1, -1, 54, -1, -1, 57, 58, -1, -1, 61, -1, -1, 64, 65, 66, 67, 68, -1, -1, 71, -1, -1, 74, 75, -1, -1, 78, -1, -1, 81, 82, 83, -1, -1, 86, -1, -1, 89, 90, -1, -1, 229, 94, 95, 96, 97, -1, -1, 100, -1, -1, 103, 104, -1, -1, 107, -1, -1, 110, 111, 112, -1, -1, 115, -1, -1, 118, 119, -1, -1, 122, -1, -1, 125, 126, 127, 128, 129, 231, 131, -1, -1, 233, 135, 136, 137, -1, -1, 140, -1, -1, 143, 144, -1, -1, 147, -1, -1, 150, 151, 152, 153, -1, -1, 156, -1, -1, 159, 160, -1, -1, 163, -1, -1, 166, 167, 168, -1, -1, 235, 172, 173, -1, -1, 237, 177, 178, 179, 180, 181, -1, -1, 184, -1, -1, 187, 188, -1, -1, 239, 192, 241, 194, 195, -1, -1, 198, -1, -1, 201, 202, 203, 204, -1, -1, 243, 208, 209, -1, -1, 212, -1, -1, 215, 216, 245, 218, -1, -1, 221, 222, -1, -1, 225, -1, -1, -1, -1, -1, -1, -1, -1, 247, 249, -1, -1, -1, -1, -1, -1, 251, 253, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((122, 59, 30, 17, 12, 9, 8, -1, -1, 11, -1, -1, 14, 220, 16, -1, -1, 23, 20, 222, 22, -1, -1, 27, 26, -1, -1, 29, -1, -1, 44, 37, 36, 35, -1, -1, 224, 41, 40, -1, -1, 43, -1, -1, 52, 49, 48, -1, -1, 51, -1, -1, 56, 55, -1, -1, 58, -1, -1, 91, 76, 69, 66, 65, -1, -1, 68, -1, -1, 73, 72, -1, -1, 75, -1, -1, 84, 81, 80, -1, -1, 83, -1, -1, 88, 87, -1, -1, 90, -1, -1, 107, 100, 97, 96, -1, -1, 99, -1, -1, 104, 103, -1, -1, 106, -1, -1, 115, 112, 111, -1, -1, 114, -1, -1, 119, 118, -1, -1, 121, -1, -1, 170, 151, 138, 133, 130, 129, -1, -1, 132, -1, -1, 137, 136, -1, -1, 226, 146, 143, 142, -1, -1, 145, -1, -1, 150, 149, -1, -1, 228, 161, 154, 230, 158, 157, -1, -1, 160, -1, -1, 169, 166, 165, -1, -1, 168, -1, -1, 232, 198, 187, 180, 177, 176, -1, -1, 179, -1, -1, 184, 183, -1, -1, 186, -1, -1, 193, 190, 234, 192, -1, -1, 197, 196, -1, -1, 236, 212, 207, 204, 203, -1, -1, 206, -1, -1, 211, 210, -1, -1, 238, 214, 240, 216, 242, 218, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 244, 246, 248, 250, -1, -1, -1, -1, -1, -1, 252, 254, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (112, 61, 32, 19, 12, 9, 8, -1, -1, 11, -1, -1, 16, 15, -1, -1, 18, -1, -1, 27, 24, 23, -1, -1, 26, -1, -1, 31, 30, -1, -1, 214, 46, 39, 36, 216, 38, -1, -1, 43, 42, -1, -1, 45, -1, -1, 54, 51, 50, -1, -1, 53, -1, -1, 58, 57, -1, -1, 60, -1, -1, 89, 76, 71, 68, 67, -1, -1, 70, -1, -1, 73, 218, 75, -1, -1, 82, 79, 220, 81, -1, -1, 86, 85, -1, -1, 88, -1, -1, 103, 98, 95, 94, -1, -1, 97, -1, -1, 100, 222, 102, -1, -1, 105, 224, 109, 108, -1, -1, 111, -1, -1, 166, 137, 126, 119, 118, 226, 228, 123, 122, -1, -1, 125, -1, -1, 130, 129, 230, 232, 134, 133, -1, -1, 136, -1, -1, 151, 146, 143, 142, -1, -1, 145, -1, -1, 150, 149, -1, -1, 234, 159, 156, 155, -1, -1, 158, -1, -1, 163, 162, -1, -1, 165, -1, -1, 192, 183, 176, 173, 172, -1, -1, 175, -1, -1, 180, 179, -1, -1, 182, -1, -1, 191, 188, 187, -1, -1, 190, -1, -1, 236, 200, 199, 196, 238, 198, -1, -1, 240, 208, 205, 204, -1, -1, 207, -1, -1, 212, 211, -1, -1, 242, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 244, 246, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 248, 250, -1, -1, 252, 254, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (124, 63, 32, 19, 12, 9, 8, -1, -1, 11, -1, -1, 16, 15, -1, -1, 18, -1, -1, 27, 24, 23, -1, -1, 26, -1, -1, 31, 30, -1, -1, 228, 48, 41, 38, 37, -1, -1, 40, -1, -1, 45, 44, -1, -1, 47, -1, -1, 56, 53, 52, -1, -1, 55, -1, -1, 60, 59, -1, -1, 62, -1, -1, 93, 80, 73, 70, 69, -1, -1, 72, -1, -1, 77, 76, -1, -1, 79, -1, -1, 88, 85, 84, -1, -1, 87, -1, -1, 92, 91, -1, -1, 230, 109, 102, 99, 98, -1, -1, 101, -1, -1, 106, 105, -1, -1, 108, -1, -1, 117, 114, 113, -1, -1, 116, -1, -1, 121, 120, -1, -1, 123, -1, -1, 176, 149, 134, 133, 130, 232, 132, -1, -1, 234, 142, 139, 138, -1, -1, 141, -1, -1, 146, 145, -1, -1, 148, -1, -1, 165, 158, 155, 154, -1, -1, 157, -1, -1, 162, 161, -1, -1, 164, -1, -1, 171, 170, 169, -1, -1, 236, 175, 174, -1, -1, 238, 200, 191, 186, 183, 182, -1, -1, 185, -1, -1, 190, 189, -1, -1, 240, 193, 242, 197, 196, -1, -1, 199, -1, -1, 214, 207, 206, 205, -1, -1, 244, 211, 210, -1, -1, 213, -1, -1, 220, 217, 246, 219, -1, -1, 224, 223, -1, -1, 226, -1, -1, -1, -1, -1, -1, -1, -1, 248, 250, -1, -1, -1, -1, -1, -1, 252, 254, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 1, 2, 3, 4, 5, 6, 6, 5, 9, 9, 4, 12, 12, 14, 14, 3, 17, 18, 18, 20, 20, 17, 23, 24, 24, 23, 27, 27, 2, 30, 31, 32, 33, 33, 32, 31, 37, 38, 38, 37, 41, 41, 30, 44, 45, 46, 46, 45, 49, 49, 44, 52, 53, 53, 52, 56, 56, 1, 59, 60, 61, 62, 63, 63, 62, 66, 66, 61, 69, 70, 70, 69, 73, 73, 60, 76, 77, 78, 78, 77, 81, 81, 76, 84, 85, 85, 84, 88, 88, 59, 91, 92, 93, 94, 94, 93, 97, 97, 92, 100, 101, 101, 100, 104, 104, 91, 107, 108, 109, 109, 108, 112, 112, 107, 115, 116, 116, 115, 119, 119, 0, 122, 123, 124, 125, 126, 127, 127, 126, 130, 130, 125, 133, 134, 134, 133, 124, 138, 139, 140, 140, 139, 143, 143, 138, 146, 147, 147, 146, 123, 151, 152, 152, 154, 155, 155, 154, 158, 158, 151, 161, 162, 163, 163, 162, 166, 166, 161, 122, 170, 171, 172, 173, 174, 174, 173, 177, 177, 172, 180, 181, 181, 180, 184, 184, 171, 187, 188, 188, 190, 190, 187, 193, 194, 194, 193, 170, 198, 199, 200, 201, 201, 200, 204, 204, 199, 207, 208, 208, 207, 198, 212, 212, 214, 214, 216, 216, 13, 13, 19, 19, 36, 36, 137, 137, 150, 150, 153, 153, 169, 169, 189, 189, 197, 197, 211, 211, 213, 213, 215, 215, 229, 229, 230, 230, 231, 231, 232, 232, 239, 239, 240, 240),
                (-1, 0, 1, 2, 3, 4, 5, 6, 6, 5, 9, 9, 4, 12, 13, 13, 12, 16, 16, 3, 19, 20, 21, 21, 20, 24, 24, 19, 27, 28, 28, 27, 2, 32, 33, 34, 34, 36, 36, 33, 39, 40, 40, 39, 43, 43, 32, 46, 47, 48, 48, 47, 51, 51, 46, 54, 55, 55, 54, 58, 58, 1, 61, 62, 63, 64, 65, 65, 64, 68, 68, 63, 71, 71, 73, 73, 62, 76, 77, 77, 79, 79, 76, 82, 83, 83, 82, 86, 86, 61, 89, 90, 91, 92, 92, 91, 95, 95, 90, 98, 98, 100, 100, 89, 103, 103, 105, 106, 106, 105, 109, 109, 0, 112, 113, 114, 115, 116, 116, 115, 119, 120, 120, 119, 123, 123, 114, 126, 127, 127, 126, 130, 131, 131, 130, 134, 134, 113, 137, 138, 139, 140, 140, 139, 143, 143, 138, 146, 147, 147, 146, 137, 151, 152, 153, 153, 152, 156, 156, 151, 159, 160, 160, 159, 163, 163, 112, 166, 167, 168, 169, 170, 170, 169, 173, 173, 168, 176, 177, 177, 176, 180, 180, 167, 183, 184, 185, 185, 184, 188, 188, 183, 166, 192, 193, 194, 194, 196, 196, 193, 192, 200, 201, 202, 202, 201, 205, 205, 200, 208, 209, 209, 208, 31, 31, 35, 35, 72, 72, 78, 78, 99, 99, 104, 104, 117, 117, 118, 118, 128, 128, 129, 129, 150, 150, 191, 191, 195, 195, 199, 199, 212, 212, 223, 223, 224, 224, 235, 235, 236, 236, 239, 239, 240, 240),
                (-1, 0, 1, 2, 3, 4, 5, 6, 6, 5, 9, 9, 4, 12, 13, 13, 12, 16, 16, 3, 19, 20, 21, 21, 20, 24, 24, 19, 27, 28, 28, 27, 2, 32, 33, 34, 35, 35, 34, 38, 38, 33, 41, 42, 42, 41, 45, 45, 32, 48, 49, 50, 50, 49, 53, 53, 48, 56, 57, 57, 56, 60, 60, 1, 63, 64, 65, 66, 67, 67, 66, 70, 70, 65, 73, 74, 74, 73, 77, 77, 64, 80, 81, 82, 82, 81, 85, 85, 80, 88, 89, 89, 88, 63, 93, 94, 95, 96, 96, 95, 99, 99, 94, 102, 103, 103, 102, 106, 106, 93, 109, 110, 111, 111, 110, 114, 114, 109, 117, 118, 118, 117, 121, 121, 0, 124, 125, 126, 127, 128, 128, 130, 130, 127, 126, 134, 135, 136, 136, 135, 139, 139, 134, 142, 143, 143, 142, 146, 146, 125, 149, 150, 151, 152, 152, 151, 155, 155, 150, 158, 159, 159, 158, 162, 162, 149, 165, 166, 167, 167, 166, 165, 171, 172, 172, 171, 124, 176, 177, 178, 179, 180, 180, 179, 183, 183, 178, 186, 187, 187, 186, 177, 191, 191, 193, 194, 194, 193, 197, 197, 176, 200, 201, 202, 203, 203, 202, 201, 207, 208, 208, 207, 211, 211, 200, 214, 215, 215, 217, 217, 214, 220, 221, 221, 220, 224, 224, 31, 31, 92, 92, 129, 129, 133, 133, 170, 170, 175, 175, 190, 190, 192, 192, 206, 206, 216, 216, 233, 233, 234, 234, 241, 241, 242, 242)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 6, 7, 7, 4, 5, 6, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 6, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 1, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 3, 4, 5, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 6, 7, 7, 5, 6, 7, 7, 6, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 4, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7),
                (0, 1, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 3, 4, 5, 6, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 6, 7, 7, 4, 5, 6, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 6, 7, 7, 4, 5, 5, 6, 7, 7, 6, 7, 7, 1, 2, 3, 4, 5, 6, 6, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 6, 5, 6, 7, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 3, 4, 5, 6, 6, 7, 7, 5, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7),
                (0, 1, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 1, 2, 3, 4, 5, 6, 6, 7, 7, 5, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 7, 7, 6, 5, 6, 7, 7, 6, 2, 3, 4, 5, 6, 7, 7, 6, 7, 7, 5, 6, 7, 7, 6, 4, 5, 5, 6, 7, 7, 6, 7, 7, 3, 4, 5, 6, 7, 7, 6, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 6, 7, 7, 5, 6, 7, 7, 6, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((7, 8, 10, 11, 15, 16, 21, 22, 25, 26, 28, 29, 34, 35, 39, 40, 42, 43, 47, 48, 50, 51, 54, 55, 57, 58, 64, 65, 67, 68, 71, 72, 74, 75, 79, 80, 82, 83, 86, 87, 89, 90, 95, 96, 98, 99, 102, 103, 105, 106, 110, 111, 113, 114, 117, 118, 120, 121, 128, 129, 131, 132, 135, 136, 141, 142, 144, 145, 148, 149, 156, 157, 159, 160, 164, 165, 167, 168, 175, 176, 178, 179, 182, 183, 185, 186, 191, 192, 195, 196, 202, 203, 205, 206, 209, 210, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 233, 234, 235, 236, 237, 238, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254),
                (7, 8, 10, 11, 14, 15, 17, 18, 22, 23, 25, 26, 29, 30, 37, 38, 41, 42, 44, 45, 49, 50, 52, 53, 56, 57, 59, 60, 66, 67, 69, 70, 74, 75, 80, 81, 84, 85, 87, 88, 93, 94, 96, 97, 101, 102, 107, 108, 110, 111, 121, 122, 124, 125, 132, 133, 135, 136, 141, 142, 144, 145, 148, 149, 154, 155, 157, 158, 161, 162, 164, 165, 171, 172, 174, 175, 178, 179, 181, 182, 186, 187, 189, 190, 197, 198, 203, 204, 206, 207, 210, 211, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 237, 238, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254),
                (7, 8, 10, 11, 14, 15, 17, 18, 22, 23, 25, 26, 29, 30, 36, 37, 39, 40, 43, 44, 46, 47, 51, 52, 54, 55, 58, 59, 61, 62, 68, 69, 71, 72, 75, 76, 78, 79, 83, 84, 86, 87, 90, 91, 97, 98, 100, 101, 104, 105, 107, 108, 112, 113, 115, 116, 119, 120, 122, 123, 131, 132, 137, 138, 140, 141, 144, 145, 147, 148, 153, 154, 156, 157, 160, 161, 163, 164, 168, 169, 173, 174, 181, 182, 184, 185, 188, 189, 195, 196, 198, 199, 204, 205, 209, 210, 212, 213, 218, 219, 222, 223, 225, 226, 227, 228, 229, 230, 231, 232, 235, 236, 237, 238, 239, 240, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((1, 1, 1, 0, 0, 1, 2, -2, 0, -2, -2, -2, 1, 1, -2, 1, -2, -2, 0, -2, 1, -2, -2, 0, 0, 2, 0, -2, -2, 0, -2, -2, 1, -2, -2, 1, 2, 1, -2, -2, -2, 0, -2, -2, 2, 1, 0, -2, -2, 2, 1, 1, -2, -2, 1, -2, -2, 0, -2, 1, -2, -2, 0, 2, 0, -2, 1, -2, -2, 1, 0, -2, -2, -2, -2, 2, 0, 1, 2, 0, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, -2, 2, 1, 0, -2, -2, -2, 0, 0, -2, -2, 0, -2, -2, 2, 0, 1, 1, -2, -2, 0, -2, -2, 0, 1, -2, -2, 1, -2, -2, 1, 0, 1, -2, -2, 1, -2, -2, 1, -2, 1, -2, -2, 2, 2, 1, 1, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 1, 0, -2, 0, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 1, 1, 1, -2, -2, -2, 1, 1, -2, -2, -2, 1, 0, 0, -2, -2, -2, 1, -2, -2, 0, 2, 2, 0, 1, 2, -2, 0, -2, -2, -2, 2, 1, -2, -2, 0, 0, -2, -2, 0, -2, -2, 1, 0, 0, -2, 1, -2, -2, 1, -2, 1, -2, -2, 0, 1, 1, -2, -2, -2, 0, -2, -2, 0, 0, -2, 2, 1, -2, 1, -2, -2, 1, 1, -2, -2, 1, -2, -2, 1, 1, 0, 2, -2, -2, 1, -2, -2, 0, 0, -2, -2, 2, -2, -2, 0, 1, 0, -2, -2, 0, -2, -2, 2, 0, -2, -2, 1, -2, -2, 1, 2, 1, 0, 1, -2, 0, -2, -2, -2, 1, -2, 0, 0, -2, -2, 1, -2, -2, 0, 1, 2, 0, -2, -2, 0, -2, -2, 2, 1, -2, -2, -2, 0, 1, -2, 0, -2, -2, 0, 1, -2, -2, -2, 1, 1, 0, -2, -2, 0, -2, 1, -2, 2, -2, -2, 0, 0, 0, 1, -2, -2, 2, -2, -2, 0, 1, -2, -2, 1, -2, -2, 1, 1, -2, 1, -2, -2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 1, 0, 1, 1, 2, 1, -2, -2, 1, -2, -2, 0, 1, -2, -2, 0, -2, -2, 0, 1, 1, -2, -2, -2, 2, 1, -2, -2, 0, -2, -2, 1, -2, 1, -2, 0, 2, -2, -2, 1, -2, -2, 1, 0, 1, 0, -2, 2, -2, -2, 0, 0, -2, -2, 2, -2, -2, 1, 1, 0, -2, -2, -2, 0, -2, 2, -2, -2, 0, 0, -2, 0, -2, 0, -2, -2, 0, 0, -2, 0, -2, -2, 1, 1, -2, -2, 2, -2, -2, 1, 1, 1, 2, 0, 1, -2, -2, 0, -2, -2, 2, 0, -2, -2, 0, -2, -2, 1, 0, -2, -2, 0, -2, -2, 0, 0, -2, 1, 1, -2, -2, 2, -2, -2, 2, 0, 0, -2, -2, -2, 2, 0, -2, -2, -2, 1, 1, -2, 1, 2, 0, -2, -2, 1, -2, -2, 1, 0, -2, -2, -2, 2, 0, 1, 0, -2, -2, -2, 2, 1, -2, -2, -2, 0, 0, -2, 1, -2, -2, -2, 1, 2, 1, 0, 0, -2, 1, 0, -2, -2, 0, -2, -2, -2, 0, 0, 0, -2, 0, -2, -2, 0, -2, 1, -2, -2, 1, -2, 0, 0, -2, -2, 0, -2, -2, 1, 1, 0, 1, 0, -2, -2, -2, 0, 1, -2, -2, -2, 1, 1, -2, 0, -2, -2, 0, 1, -2, -2, 0, -2, -2, 0, 1, 0, -2, -2, 0, -2, 0, -2, -2, 1, -2, 1, -2, -2, 1, 1, -2, 1, 2, 1, 0, -2, -2, 1, -2, -2, 0, -2, -2, 0, 1, 2, -2, -2, 2, -2, -2, 1, -2, 2, -2, -2, 1, -2, 0, 0, 2, -2, 0, -2, -2, 1, 0, -2, -2, 2, -2, -2, 0, 1, 1, -2, -2, 0, -2, -2, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 1, 2, 0, 1, 0, -2, -2, -2, 0, 0, -2, -2, 0, 1, -2, -2, -2, 1, 0, -2, 0, 1, -2, -2, -2, 0, -2, 1, -2, 1, -2, -2, 0, 2, 1, 1, 0, -2, -2, 1, -2, -2, 1, 0, -2, -2, 0, -2, -2, 1, 1, 1, -2, -2, -2, 1, 0, -2, -2, -2, 2, 1, 1, -2, 0, -2, -2, 1, -2, 1, -2, -2, 0, 0, 0, -2, -2, 1, -2, -2, 1, -2, 1, -2, -2, 1, 2, 1, 1, 1, 1, -2, -2, -2, 0, 1, -2, -2, -2, 1, -2, 0, 1, -2, -2, 0, -2, -2, 0, 0, 1, 1, -2, -2, -2, 1, 1, -2, -2, 0, -2, -2, 1, 1, -2, 1, -2, -2, 2, 0, -2, -2, 1, -2, -2, 2, 1, 0, 1, -2, 1, -2, -2, -2, 1, -2, 0, 1, -2, -2, -2, 0, 2, 1, 1, -2, -2, 0, -2, -2, 0, -2, 0, -2, -2, 0, 1, 0, -2, -2, 2, -2, -2, -2, 2, 2, 1, 1, 0, 0, -2, 1, -2, -2, -2, 1, 0, -2, -2, 0, 0, -2, -2, 0, -2, -2, 0, 0, -2, 1, 0, -2, -2, 0, -2, -2, 1, 0, 0, -2, -2, 0, -2, -2, 0, -2, -2, 0, 1, 2, 1, 1, -2, -2, 1, -2, -2, 0, 1, -2, -2, 0, -2, -2, 2, 1, 1, -2, -2, -2, 0, 1, -2, -2, 0, -2, -2, 1, 2, 1, 1, -2, -2, 1, -2, -2, 0, 1, -2, -2, -2, 2, 0, 1, -2, -2, 0, -2, -2, 0, 0, -2, -2, 0, -2, -2, 1, 0, 1, 2, 1, 1, -2, -2, 0, -2, -2, 1, 1, -2, -2, 1, -2, -2, 2, 0, 0, -2, -2, -2, 0, 1, -2, -2, 0, -2, -2, 1, 1, -2, 1, -2, -2, 1, -2, 1, 1, -2, -2, 0, -2, -2, 1, -2, 2, 0, 1, 0, -2, -2, -2, 0, 0, -2, -2, -2, 0, 1, 1, -2, -2, 0, -2, -2, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((2256, 1224, 926, 3683, 1140, 123, 139, -256, 534, -256, -256, -256, 402, 255, -256, 317, -256, -256, 2546, -256, 483, -256, -256, 5760, 5391, 134, 3829, -256, -256, 4956, -256, -256, 492, -256, -256, 923, 109, 899, -256, -256, -256, 12107, -256, -256, 134, 930, 34052, -256, -256, 92, 936, 936, -256, -256, 958, -256, -256, 8906, -256, 1033, -256, -256, 8147, 164, 6894, -256, 1086, -256, -256, 1063, 5666, -256, -256, -256, -256, 109, 22954, 1477, 92, 15944, 15231, -256, -256, 17972, -256, -256, 15350, 1287, -256, -256, -256, 92, 1617, 20460, -256, -256, -256, 20675, 17777, -256, -256, 21164, -256, -256, 92, 31945, 1788, 1680, -256, -256, 29420, -256, -256, 36490, 2113, -256, -256, 2228, -256, -256, 2211, 24096, 1870, -256, -256, 2099, -256, -256, 2211, -256, 2235, -256, -256, 164, 134, 1877, 1224, -256, 15155, -256, -256, 26887, 1975, -256, -256, 28131, -256, -256, 1504, 11389, -256, 12402, -256, -256, 21845, 1811, -256, -256, 2134, -256, -256, 19178, 1776, 1763, 1549, -256, -256, -256, 2028, 2018, -256, -256, -256, 2207, 20589, 20532, -256, -256, -256, 2208, -256, -256, 44659, 134, 109, 40835, 2443, 92, -256, 35190, -256, -256, -256, 92, 2351, -256, -256, 41066, 40967, -256, -256, 43777, -256, -256, 2689, 35929, 31990, -256, 2408, -256, -256, 2603, -256, 2616, -256, -256, 44116, 2715, 2713, -256, -256, -256, 44578, -256, -256, 33104, 24682, -256, 164, 2328, -256, 2582, -256, -256, 2577, 2463, -256, -256, 2740, -256, -256, 3036, 2805, 33359, 164, -256, -256, 2669, -256, -256, 37394, 33257, -256, -256, 164, -256, -256, 43199, 3127, 36810, -256, -256, 40846, -256, -256, 164, 43328, -256, -256, 3496, -256, -256, 3069, 92, 2741, 52378, 2440, -256, 48583, -256, -256, -256, 2742, -256, 62717, 58824, -256, -256, 3033, -256, -256, 53073, 2841, 109, 46170, -256, -256, 48676, -256, -256, 134, 2985, -256, -256, -256, 55072, 2822, -256, 55034, -256, -256, 57529, 2910, -256, -256, -256, 3073, 3071, 53881, -256, -256, 50157, -256, 3072, -256, 101, -256, -256, 71782, 53761, 48564, 3116, -256, -256, 134, -256, -256, 66328, 3416, -256, -256, 3392, -256, -256, 3644, 3249, -256, 3249, -256, -256, 86368, 3662, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256),
                (134, 2363, 1635, 11325, 713, 330, 92, 262, -256, -256, 190, -256, -256, 3667, 397, -256, -256, 4916, -256, -256, 7108, 855, 849, -256, -256, -256, 92, 1023, -256, -256, 7441, -256, -256, 1208, -256, 1208, -256, 15488, 109, -256, -256, 1444, -256, -256, 1912, 23742, 1645, 18703, -256, 92, -256, -256, 21212, 17659, -256, -256, 92, -256, -256, 1870, 1656, 24293, -256, -256, -256, 26183, -256, 92, -256, -256, 29641, 24683, -256, 25458, -256, 26890, -256, -256, 33820, 30674, -256, 33403, -256, -256, 2356, 2222, -256, -256, 109, -256, -256, 3003, 2745, 2719, 92, 46165, 2416, -256, -256, 52057, -256, -256, 109, 42902, -256, -256, 38238, -256, -256, 2729, 34377, -256, -256, 46563, -256, -256, 52830, 44142, -256, 2875, 2873, -256, -256, 109, -256, -256, 92, 62166, 57097, -256, -256, -256, 109, 55680, -256, -256, -256, 3478, 3004, -256, 3460, 92, 75827, -256, -256, 3220, -256, -256, 3476, 67978, -256, -256, -256, 109, 86994, 3619, 74990, -256, -256, -256, 92, 3500, -256, -256, -256, 65327, 63419, -256, 3593, -256, -256, -256, 2276, 164, 1086, 6498, 1239, -256, 528, 1915, -256, -256, 4919, -256, -256, -256, 16623, 10445, 8972, -256, 9011, -256, -256, 10493, -256, 1552, -256, -256, 1820, -256, 21789, 20348, -256, -256, 24937, -256, -256, 1730, 731, 2501, 329, 664, -256, -256, -256, 2758, 421, -256, -256, -256, 732, 732, -256, 75985, -256, -256, 8559, 1063, -256, -256, 11649, -256, -256, 19162, 1735, 14883, -256, -256, 17135, -256, 17728, -256, -256, 2203, -256, 2204, -256, -256, 2948, 2276, -256, 2289, 164, 2286, 25691, -256, -256, 2288, -256, -256, 30065, -256, -256, 32109, 2434, 164, -256, -256, 164, -256, -256, 2734, -256, 164, -256, -256, 2948, -256, 43471, 39788, 164, -256, 37491, -256, -256, 3224, 42073, -256, -256, 164, -256, -256, 49668, 3341, 3172, -256, -256, 46098, -256, -256, 53900, 53842, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256),
                (2194, 109, 993, 92, 5255, 551, 1247, -256, -256, -256, 6279, 6202, -256, -256, 9658, 902, -256, -256, -256, 677, 1159, -256, 3857, 489, -256, -256, -256, 6284, -256, 955, -256, 956, -256, -256, 21727, 92, 1372, 1021, 8445, -256, -256, 1368, -256, -256, 1499, 18026, -256, -256, 21611, -256, -256, 1465, 1460, 1402, -256, -256, -256, 1651, 18537, -256, -256, -256, 92, 1777, 1683, -256, 24428, -256, -256, 1778, -256, 2000, -256, -256, 26777, 25774, 25536, -256, -256, 1456, -256, -256, 2029, -256, 2030, -256, -256, 1558, 134, 832, 441, 267, 267, -256, -256, -256, 4468, 531, -256, -256, -256, 832, -256, 11453, 1089, -256, -256, 13769, -256, -256, 6483, 2427, 224, 163, -256, -256, -256, 722, 659, -256, -256, 6381, -256, -256, 1300, 1136, -256, 1136, -256, -256, 164, 13294, -256, -256, 1369, -256, -256, 134, 1812, 18026, 1657, -256, 1664, -256, -256, -256, 1813, -256, 27445, 1833, -256, -256, -256, 19099, 164, 1647, 1643, -256, -256, 17735, -256, -256, 14316, -256, 16672, -256, -256, 21845, 2044, 20552, -256, -256, 164, -256, -256, -256, 134, 92, 2775, 2228, 39065, 35425, -256, 2221, -256, -256, -256, 2251, 42348, -256, -256, 49934, 42253, -256, -256, 52063, -256, -256, 76491, 58903, -256, 3079, 62717, -256, -256, 72843, -256, -256, 3789, 84613, 77963, -256, -256, 89603, -256, -256, 116240, -256, -256, 53801, 2691, 109, 2680, 2641, -256, -256, 2680, -256, -256, 34761, 2209, -256, -256, 38238, -256, -256, 109, 2831, 2804, -256, -256, -256, 44410, 2715, -256, -256, 44533, -256, -256, 3303, 109, 3095, 2827, -256, -256, 3096, -256, -256, 58795, 3175, -256, -256, -256, 109, 71915, 3496, -256, -256, 76917, -256, -256, 64052, 59511, -256, -256, 66388, -256, -256, 2937, 28355, 2239, 164, 2227, 2200, -256, -256, 14059, -256, -256, 2203, 2199, -256, -256, 2227, -256, -256, 164, 28301, 26782, -256, -256, -256, 27969, 2495, -256, -256, 28277, -256, -256, 2667, 2648, -256, 2649, -256, -256, 2667, -256, 2668, 2668, -256, -256, 38318, -256, -256, 2938, -256, 164, 45934, 3129, 40842, -256, -256, -256, 55320, 55254, -256, -256, -256, 42312, 3036, 3035, -256, -256, 40339, -256, -256, 3438, -256, 3439, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256, -256)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((38, 41, 42, 42, 13, 1, 4, 0, 5, 0, 43, 0, 19, 35, 43, 22, 0, 29, 1, 0, 2, 21, 0, 43, 35, 35, 34, 43, 32, 38, 35, 41, 11, 43, 0, 43, 43, 43, 43, 42, 43, 42, 0, 43, 41, 41, 32, 0, 43, 41, 41, 38, 43, 0, 41, 43, 41, 41, 0, 43, 43, 43, 41, 4, 4, 0, 18, 43, 0, 3, 12, 0, 43, 0, 43, 39, 39, 5, 15, 14, 1, 0, 11, 39, 28, 43, 16, 2, 8, 0, 43, 1, 0, 2, 0, 43, 0, 2, 0, 0, 3, 19, 43, 13, 42, 42, 24, 42, 43, 36, 5, 0, 16, 42, 36, 42, 0, 43, 43, 42, 42, 42, 26, 43, 0, 43, 43, 42, 40, 0, 41, 42, 39, 40, 39, 39, 40, 0, 40, 1, 42, 38, 0, 1, 0, 43, 36, 43, 40, 41, 0, 43, 32, 43, 39, 4, 10, 0, 43, 43, 42, 40, 7, 14, 14, 17, 7, 43, 1, 1, 1, 43, 0, 43, 43, 39, 43, 0, 43, 42, 0, 43, 34, 4, 2, 1, 0, 1, 0, 1, 0, 21, 0, 7, 2, 43, 0, 11, 34, 43, 28, 9, 11, 0, 3, 9, 1, 0, 12, 34, 0, 40, 43, 34, 0, 36, 0, 0, 3, 0, 43, 0, 28, 43, 0, 7, 2, 0, 8, 5, 43, 3, 14, 0, 13, 39, 43, 30, 2, 17, 0, 23, 37, 41, 28, 14, 43, 41, 43, 38, 27, 13, 43, 11, 39, 32, 43, 5, 2, 9, 0, 14, 1, 0, 5, 22, 16, 43, 7, 27, 43, 0, 41, 42, 41, 42, 23, 43, 8, 0, 12, 43, 39, 0, 39, 6, 2, 17, 43, 43, 42, 42, 38, 42, 40, 28, 43, 42, 42, 43, 27, 9, 11, 0, 43, 43, 42, 43, 39, 43, 0, 43, 42, 43, 40, 43, 40, 30, 38, 0, 43, 21, 0, 36, 43, 21, 0, 43, 40, 22, 14, 9, 34, 8, 18, 0, 37, 26, 24, 26, 19, 31, 35, 26, 42, 42, 43, 42, 34, 42, 41, 20, 0, 28, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0),
                (38, 37, 40, 41, 16, 33, 36, 35, 37, 28, 37, 34, 40, 29, 1, 5, 0, 42, 38, 43, 4, 0, 1, 0, 43, 0, 11, 12, 40, 0, 10, 43, 9, 42, 43, 42, 0, 42, 7, 3, 13, 43, 43, 42, 37, 38, 2, 14, 0, 36, 0, 43, 2, 0, 0, 3, 13, 0, 26, 42, 43, 42, 0, 43, 43, 42, 0, 42, 42, 43, 37, 1, 0, 9, 43, 8, 3, 10, 42, 26, 43, 23, 25, 7, 43, 43, 43, 42, 41, 40, 43, 32, 34, 35, 35, 34, 0, 2, 0, 42, 26, 43, 35, 35, 1, 43, 35, 2, 43, 38, 42, 0, 43, 37, 0, 43, 33, 2, 0, 14, 20, 19, 43, 7, 0, 28, 42, 41, 15, 6, 23, 43, 43, 43, 38, 43, 43, 30, 31, 0, 31, 31, 29, 1, 42, 32, 33, 31, 35, 34, 0, 42, 43, 28, 27, 3, 3, 0, 27, 0, 42, 42, 40, 42, 43, 30, 0, 0, 21, 0, 43, 43, 39, 41, 41, 42, 15, 0, 21, 39, 28, 43, 6, 0, 16, 43, 40, 4, 1, 0, 5, 43, 2, 14, 43, 12, 35, 2, 42, 43, 42, 4, 0, 14, 42, 30, 43, 41, 42, 42, 9, 21, 0, 43, 0, 43, 32, 43, 0, 43, 41, 9, 0, 14, 0, 43, 41, 4, 9, 0, 42, 31, 43, 39, 1, 7, 0, 43, 0, 0, 4, 43, 0, 43, 43, 42, 0, 43, 36, 37, 0, 37, 34, 33, 37, 0, 43, 19, 24, 0, 35, 0, 43, 37, 3, 9, 4, 13, 1, 1, 2, 42, 43, 42, 41, 42, 35, 0, 35, 1, 0, 0, 1, 0, 7, 15, 28, 19, 38, 3, 0, 9, 42, 28, 37, 43, 28, 13, 4, 17, 43, 39, 39, 14, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
                (38, 41, 40, 42, 42, 15, 30, 0, 43, 0, 43, 30, 43, 0, 43, 41, 43, 0, 43, 42, 42, 0, 43, 31, 43, 0, 43, 42, 0, 43, 43, 42, 0, 43, 39, 6, 6, 15, 30, 0, 43, 13, 13, 43, 1, 6, 0, 43, 0, 0, 43, 7, 15, 15, 15, 7, 43, 1, 5, 1, 43, 0, 42, 42, 43, 43, 42, 0, 43, 41, 0, 41, 41, 40, 42, 30, 32, 30, 40, 13, 43, 5, 43, 43, 42, 0, 42, 41, 42, 42, 42, 42, 42, 42, 0, 43, 42, 2, 6, 0, 43, 41, 0, 41, 7, 15, 0, 43, 30, 43, 42, 13, 1, 9, 5, 43, 0, 21, 41, 42, 32, 1, 1, 12, 43, 43, 43, 42, 0, 42, 42, 42, 5, 43, 42, 40, 42, 39, 39, 40, 1, 0, 1, 43, 0, 43, 38, 0, 39, 3, 21, 2, 43, 40, 3, 3, 12, 8, 43, 0, 0, 9, 3, 0, 16, 11, 23, 43, 34, 40, 38, 43, 9, 0, 28, 43, 35, 33, 32, 35, 40, 4, 0, 21, 43, 0, 43, 34, 27, 0, 43, 35, 2, 0, 14, 43, 33, 43, 30, 3, 0, 11, 32, 17, 41, 2, 0, 11, 42, 42, 28, 43, 26, 43, 41, 43, 18, 0, 43, 34, 6, 14, 11, 11, 12, 1, 32, 43, 21, 16, 2, 10, 1, 41, 36, 43, 2, 1, 4, 1, 14, 0, 3, 0, 3, 0, 13, 43, 12, 42, 42, 42, 43, 43, 42, 41, 0, 41, 42, 36, 41, 7, 43, 39, 38, 2, 3, 0, 42, 28, 43, 41, 9, 2, 14, 42, 30, 43, 36, 38, 2, 8, 8, 2, 9, 0, 34, 0, 43, 8, 21, 0, 43, 6, 0, 14, 1, 0, 0, 0, 5, 43, 2, 1, 3, 0, 34, 43, 0, 42, 43, 43, 42, 0, 43, 41, 0, 41, 34, 43, 0, 41, 16, 43, 35, 0, 35, 35, 2, 5, 0, 40, 0, 42, 34, 34, 0, 43, 35, 2, 9, 6, 43, 1, 0, 14, 42, 43, 42, 0, 42, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 43, 43, 0, 0, 43, 43, 43, 43, 43, 43, 0, 0, 43, 43, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 43, 43, 43, 43, 0, 0, 0, 0, 43, 43, 43, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 3, 4, 5, 6, 7, 355, 9, -1, -1, 357, 13, 14, 359, 16, -1, -1, 19, 361, 21, -1, -1, 24, 25, 26, 27, -1, -1, 30, -1, -1, 33, 363, 365, 36, 37, 38, -1, -1, 367, 42, 369, 371, 45, 46, 47, 373, 375, 50, 51, 52, -1, -1, 55, -1, -1, 58, 377, 60, -1, -1, 63, 64, 65, 379, 67, -1, -1, 70, 71, -1, -1, 381, 383, 76, 77, 78, 79, 80, 81, -1, -1, 84, -1, -1, 87, 88, -1, -1, 385, 92, 93, 94, -1, -1, 387, 98, 99, -1, -1, 102, -1, -1, 105, 106, 107, 108, -1, -1, 111, -1, -1, 114, 115, -1, -1, 118, -1, -1, 121, 122, 123, -1, -1, 126, -1, -1, 129, 389, 131, -1, -1, 134, 135, 136, 137, 391, 139, -1, -1, 142, 143, -1, -1, 146, -1, -1, 149, 150, 393, 152, -1, -1, 155, 156, -1, -1, 159, -1, -1, 162, 163, 164, 165, -1, -1, 395, 169, 170, -1, -1, 397, 174, 175, 176, -1, -1, 399, 180, 401, 403, 183, 184, 185, 186, 187, 188, 405, 190, -1, -1, 407, 194, 195, 409, 411, 198, 199, -1, -1, 202, -1, -1, 205, 206, 207, 413, 209, -1, -1, 212, 415, 214, -1, -1, 217, 218, 219, -1, -1, 417, 223, 419, 421, 226, 227, 423, 229, 230, 425, 232, -1, -1, 235, 236, -1, -1, 239, -1, -1, 242, 243, 244, 245, -1, -1, 248, -1, -1, 251, 252, -1, -1, 255, -1, -1, 258, 259, 260, -1, -1, 263, -1, -1, 266, 267, -1, -1, 270, -1, -1, 273, 274, 275, 276, 277, 427, 279, -1, -1, 429, 283, 431, 285, 286, -1, -1, 289, -1, -1, 292, 293, 294, 295, -1, -1, 298, -1, -1, 301, 302, -1, -1, 433, 306, 307, 435, 309, -1, -1, 312, 313, -1, -1, 437, 317, 318, 319, 439, 441, 322, 443, 324, 445, 326, -1, -1, 329, 330, 331, 332, -1, -1, 335, -1, -1, 338, 339, -1, -1, 342, -1, -1, 345, 346, 447, 348, -1, -1, 351, 352, -1, -1, 449, -1, -1, 451, 453, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 455, 457, 459, 461, -1, -1, -1, -1, -1, -1, 463, 465, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 467, 469, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 471, 473, -1, -1, -1, -1, 475, 477, 479, 481, -1, -1, -1, -1, -1, -1, 483, 485, 487, 489, 491, 493, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 495, 497, 499, 501, -1, -1, -1, -1, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, 7, 8, -1, -1, 11, -1, -1, 14, 15, -1, -1, 18, -1, -1, 21, 22, 23, -1, -1, 305, 27, 28, -1, -1, 31, -1, -1, 34, 307, 36, 309, 38, 39, -1, -1, 42, -1, -1, 45, 46, 47, 48, 311, 50, -1, -1, 53, 54, -1, -1, 57, -1, -1, 60, 61, 62, -1, -1, 313, 66, 315, 68, -1, -1, 71, 72, 317, 74, 319, 76, -1, -1, 79, 80, 321, 82, -1, -1, 85, 86, -1, -1, 89, -1, -1, 92, 93, 94, 95, 96, 97, -1, -1, 100, -1, -1, 103, 104, -1, -1, 107, -1, -1, 110, 111, 323, 325, 114, 327, 329, 117, 118, 331, 120, 121, -1, -1, 124, -1, -1, 127, 128, 129, -1, -1, 333, 133, 134, -1, -1, 335, 138, 139, 337, 141, 142, 143, -1, -1, 146, -1, -1, 149, 150, -1, -1, 339, 154, 155, 156, 157, -1, -1, 341, 161, 162, -1, -1, 343, 166, 167, 345, 169, -1, -1, 347, 173, 174, 175, 176, 177, 349, 179, 180, -1, -1, 183, -1, -1, 351, 187, 188, 189, 353, 191, -1, -1, 194, 355, 196, -1, -1, 199, 357, 201, 202, -1, -1, 205, -1, -1, 208, 209, 210, 211, 212, -1, -1, 359, 216, 217, -1, -1, 361, 221, 222, 363, 224, -1, -1, 227, 228, -1, -1, 231, -1, -1, 234, 235, 236, 365, 367, 239, 369, 241, -1, -1, 244, 371, 246, 373, 375, 249, 250, 377, 252, 253, 254, 255, -1, -1, 258, -1, -1, 261, 379, 381, 264, 265, 266, -1, -1, 269, -1, -1, 272, 383, 274, -1, -1, 277, 385, 279, 280, 281, 387, 283, -1, -1, 286, 287, -1, -1, 290, -1, -1, 293, 294, 295, -1, -1, 298, -1, -1, 301, 302, -1, -1, 389, -1, -1, 391, 393, 395, 397, -1, -1, -1, -1, -1, -1, 399, 401, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 403, 405, -1, -1, -1, -1, 407, 409, -1, -1, -1, -1, -1, -1, -1, -1, 411, 413, 415, 417, 419, 421, -1, -1, -1, -1, 423, 425, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 427, 429, -1, -1, -1, -1, 431, 433, -1, -1, -1, -1, -1, -1, 435, 437, -1, -1, -1, -1, 439, 441, 443, 445, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 447, 449, 451, 453, -1, -1, -1, -1, -1, -1, -1, -1, 455, 457, 459, 461, -1, -1, -1, -1, -1, -1, -1, -1, 463, 465, 467, 469, 471, 473, 475, 477, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 2, 3, 4, 5, 6, 7, 351, 353, 355, 11, 12, 357, 359, 15, 16, -1, -1, 361, 20, 21, 363, 23, 24, -1, -1, 365, 28, 367, 30, 369, 32, -1, -1, 35, 36, 37, 38, 39, -1, -1, 42, -1, -1, 45, 46, -1, -1, 49, -1, -1, 52, 53, 54, -1, -1, 371, 58, 59, -1, -1, 373, 63, 64, 65, 375, 67, -1, -1, 70, 377, 72, -1, -1, 75, 76, 77, -1, -1, 80, -1, -1, 83, 379, 85, -1, -1, 88, 89, 90, 91, 92, 93, -1, -1, 381, 97, 98, -1, -1, 383, 102, 385, 104, 105, -1, -1, 108, -1, -1, 111, 112, 113, 114, -1, -1, 387, 118, 119, -1, -1, 122, -1, -1, 125, 126, 389, 128, -1, -1, 131, 132, -1, -1, 135, -1, -1, 138, 139, 140, 141, 391, 143, -1, -1, 393, 147, 395, 149, 150, -1, -1, 397, 154, 155, 156, 157, -1, -1, 160, -1, -1, 163, 399, 165, -1, -1, 168, 169, 170, -1, -1, 173, -1, -1, 401, 177, 178, 179, 180, 181, 182, 403, 184, -1, -1, 405, 188, 189, 407, 409, 192, 193, -1, -1, 196, -1, -1, 199, 200, 411, 202, 203, -1, -1, 206, -1, -1, 209, 210, 211, -1, -1, 214, -1, -1, 217, 413, 415, 220, 221, 222, 223, 224, -1, -1, 227, -1, -1, 230, 231, -1, -1, 234, -1, -1, 237, 238, 239, -1, -1, 417, 243, 244, -1, -1, 247, -1, -1, 250, 251, 252, 253, -1, -1, 256, -1, -1, 259, 260, -1, -1, 419, 264, 265, 266, -1, -1, 269, -1, -1, 272, 273, -1, -1, 276, -1, -1, 279, 280, 281, 282, 283, 284, -1, -1, 287, -1, -1, 290, 291, -1, -1, 294, -1, -1, 297, 298, 299, -1, -1, 421, 303, 304, -1, -1, 307, -1, -1, 310, 311, 423, 313, 425, 427, 316, 429, 318, 319, -1, -1, 322, -1, -1, 325, 431, 327, 328, 329, 330, -1, -1, 433, 334, 335, -1, -1, 435, 339, 340, 341, -1, -1, 344, -1, -1, 347, 437, 349, -1, -1, -1, -1, -1, -1, 439, 441, -1, -1, -1, -1, -1, -1, 443, 445, -1, -1, 447, 449, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 451, 453, -1, -1, -1, -1, -1, -1, 455, 457, 459, 461, -1, -1, -1, -1, 463, 465, -1, -1, 467, 469, -1, -1, -1, -1, 471, 473, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 475, 477, -1, -1, -1, -1, 479, 481, 483, 485, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((182, 75, 44, 23, 12, 11, 8, 356, 10, -1, -1, 358, 18, 15, 360, 17, -1, -1, 20, 362, 22, -1, -1, 35, 32, 29, 28, -1, -1, 31, -1, -1, 34, 364, 366, 41, 40, 39, -1, -1, 368, 43, 370, 372, 62, 49, 48, 374, 376, 57, 54, 53, -1, -1, 56, -1, -1, 59, 378, 61, -1, -1, 74, 69, 66, 380, 68, -1, -1, 73, 72, -1, -1, 382, 384, 133, 104, 91, 86, 83, 82, -1, -1, 85, -1, -1, 90, 89, -1, -1, 386, 97, 96, 95, -1, -1, 388, 101, 100, -1, -1, 103, -1, -1, 120, 113, 110, 109, -1, -1, 112, -1, -1, 117, 116, -1, -1, 119, -1, -1, 128, 125, 124, -1, -1, 127, -1, -1, 130, 390, 132, -1, -1, 161, 148, 141, 138, 392, 140, -1, -1, 145, 144, -1, -1, 147, -1, -1, 154, 151, 394, 153, -1, -1, 158, 157, -1, -1, 160, -1, -1, 173, 168, 167, 166, -1, -1, 396, 172, 171, -1, -1, 398, 179, 178, 177, -1, -1, 400, 181, 402, 404, 272, 225, 204, 193, 192, 189, 406, 191, -1, -1, 408, 197, 196, 410, 412, 201, 200, -1, -1, 203, -1, -1, 216, 211, 208, 414, 210, -1, -1, 213, 416, 215, -1, -1, 222, 221, 220, -1, -1, 418, 224, 420, 422, 241, 228, 424, 234, 231, 426, 233, -1, -1, 238, 237, -1, -1, 240, -1, -1, 257, 250, 247, 246, -1, -1, 249, -1, -1, 254, 253, -1, -1, 256, -1, -1, 265, 262, 261, -1, -1, 264, -1, -1, 269, 268, -1, -1, 271, -1, -1, 316, 291, 282, 281, 278, 428, 280, -1, -1, 430, 284, 432, 288, 287, -1, -1, 290, -1, -1, 305, 300, 297, 296, -1, -1, 299, -1, -1, 304, 303, -1, -1, 434, 311, 308, 436, 310, -1, -1, 315, 314, -1, -1, 438, 328, 321, 320, 440, 442, 323, 444, 325, 446, 327, -1, -1, 344, 337, 334, 333, -1, -1, 336, -1, -1, 341, 340, -1, -1, 343, -1, -1, 350, 347, 448, 349, -1, -1, 354, 353, -1, -1, 450, -1, -1, 452, 454, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 456, 458, 460, 462, -1, -1, -1, -1, -1, -1, 464, 466, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 468, 470, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 472, 474, -1, -1, -1, -1, 476, 478, 480, 482, -1, -1, -1, -1, -1, -1, 484, 486, 488, 490, 492, 494, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 496, 498, 500, 502, -1, -1, -1, -1, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (172, 91, 44, 33, 20, 13, 10, 9, -1, -1, 12, -1, -1, 17, 16, -1, -1, 19, -1, -1, 26, 25, 24, -1, -1, 306, 30, 29, -1, -1, 32, -1, -1, 35, 308, 37, 310, 41, 40, -1, -1, 43, -1, -1, 70, 59, 52, 49, 312, 51, -1, -1, 56, 55, -1, -1, 58, -1, -1, 65, 64, 63, -1, -1, 314, 67, 316, 69, -1, -1, 78, 73, 318, 75, 320, 77, -1, -1, 84, 81, 322, 83, -1, -1, 88, 87, -1, -1, 90, -1, -1, 137, 116, 109, 102, 99, 98, -1, -1, 101, -1, -1, 106, 105, -1, -1, 108, -1, -1, 113, 112, 324, 326, 115, 328, 330, 126, 119, 332, 123, 122, -1, -1, 125, -1, -1, 132, 131, 130, -1, -1, 334, 136, 135, -1, -1, 336, 153, 140, 338, 148, 145, 144, -1, -1, 147, -1, -1, 152, 151, -1, -1, 340, 165, 160, 159, 158, -1, -1, 342, 164, 163, -1, -1, 344, 171, 168, 346, 170, -1, -1, 348, 248, 207, 186, 185, 178, 350, 182, 181, -1, -1, 184, -1, -1, 352, 198, 193, 190, 354, 192, -1, -1, 195, 356, 197, -1, -1, 200, 358, 204, 203, -1, -1, 206, -1, -1, 233, 220, 215, 214, 213, -1, -1, 360, 219, 218, -1, -1, 362, 226, 223, 364, 225, -1, -1, 230, 229, -1, -1, 232, -1, -1, 243, 238, 237, 366, 368, 240, 370, 242, -1, -1, 245, 372, 247, 374, 376, 276, 251, 378, 263, 260, 257, 256, -1, -1, 259, -1, -1, 262, 380, 382, 271, 268, 267, -1, -1, 270, -1, -1, 273, 384, 275, -1, -1, 278, 386, 292, 285, 282, 388, 284, -1, -1, 289, 288, -1, -1, 291, -1, -1, 300, 297, 296, -1, -1, 299, -1, -1, 304, 303, -1, -1, 390, -1, -1, 392, 394, 396, 398, -1, -1, -1, -1, -1, -1, 400, 402, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 404, 406, -1, -1, -1, -1, 408, 410, -1, -1, -1, -1, -1, -1, -1, -1, 412, 414, 416, 418, 420, 422, -1, -1, -1, -1, 424, 426, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 428, 430, -1, -1, -1, -1, 432, 434, -1, -1, -1, -1, -1, -1, 436, 438, -1, -1, -1, -1, 440, 442, 444, 446, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 448, 450, 452, 454, -1, -1, -1, -1, -1, -1, -1, -1, 456, 458, 460, 462, -1, -1, -1, -1, -1, -1, -1, -1, 464, 466, 468, 470, 472, 474, 476, 478, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (176, 87, 34, 19, 10, 9, 8, 352, 354, 356, 14, 13, 358, 360, 18, 17, -1, -1, 362, 27, 22, 364, 26, 25, -1, -1, 366, 29, 368, 31, 370, 33, -1, -1, 62, 51, 44, 41, 40, -1, -1, 43, -1, -1, 48, 47, -1, -1, 50, -1, -1, 57, 56, 55, -1, -1, 372, 61, 60, -1, -1, 374, 74, 69, 66, 376, 68, -1, -1, 71, 378, 73, -1, -1, 82, 79, 78, -1, -1, 81, -1, -1, 84, 380, 86, -1, -1, 137, 110, 101, 96, 95, 94, -1, -1, 382, 100, 99, -1, -1, 384, 103, 386, 107, 106, -1, -1, 109, -1, -1, 124, 117, 116, 115, -1, -1, 388, 121, 120, -1, -1, 123, -1, -1, 130, 127, 390, 129, -1, -1, 134, 133, -1, -1, 136, -1, -1, 153, 146, 145, 142, 392, 144, -1, -1, 394, 148, 396, 152, 151, -1, -1, 398, 167, 162, 159, 158, -1, -1, 161, -1, -1, 164, 400, 166, -1, -1, 175, 172, 171, -1, -1, 174, -1, -1, 402, 278, 219, 198, 187, 186, 183, 404, 185, -1, -1, 406, 191, 190, 408, 410, 195, 194, -1, -1, 197, -1, -1, 208, 201, 412, 205, 204, -1, -1, 207, -1, -1, 216, 213, 212, -1, -1, 215, -1, -1, 218, 414, 416, 249, 236, 229, 226, 225, -1, -1, 228, -1, -1, 233, 232, -1, -1, 235, -1, -1, 242, 241, 240, -1, -1, 418, 246, 245, -1, -1, 248, -1, -1, 263, 258, 255, 254, -1, -1, 257, -1, -1, 262, 261, -1, -1, 420, 271, 268, 267, -1, -1, 270, -1, -1, 275, 274, -1, -1, 277, -1, -1, 324, 309, 296, 289, 286, 285, -1, -1, 288, -1, -1, 293, 292, -1, -1, 295, -1, -1, 302, 301, 300, -1, -1, 422, 306, 305, -1, -1, 308, -1, -1, 315, 312, 424, 314, 426, 428, 317, 430, 321, 320, -1, -1, 323, -1, -1, 326, 432, 338, 333, 332, 331, -1, -1, 434, 337, 336, -1, -1, 436, 346, 343, 342, -1, -1, 345, -1, -1, 348, 438, 350, -1, -1, -1, -1, -1, -1, 440, 442, -1, -1, -1, -1, -1, -1, 444, 446, -1, -1, 448, 450, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 452, 454, -1, -1, -1, -1, -1, -1, 456, 458, 460, 462, -1, -1, -1, -1, 464, 466, -1, -1, 468, 470, -1, -1, -1, -1, 472, 474, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 476, 478, -1, -1, -1, -1, 480, 482, 484, 486, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 1, 2, 3, 4, 5, 6, 6, 8, 8, 5, 4, 12, 13, 13, 15, 15, 12, 18, 18, 20, 20, 3, 23, 24, 25, 26, 26, 25, 29, 29, 24, 32, 32, 23, 35, 36, 37, 37, 36, 35, 41, 41, 2, 44, 45, 46, 46, 45, 49, 50, 51, 51, 50, 54, 54, 49, 57, 57, 59, 59, 44, 62, 63, 64, 64, 66, 66, 63, 69, 70, 70, 69, 62, 1, 75, 76, 77, 78, 79, 80, 80, 79, 83, 83, 78, 86, 87, 87, 86, 77, 91, 92, 93, 93, 92, 91, 97, 98, 98, 97, 101, 101, 76, 104, 105, 106, 107, 107, 106, 110, 110, 105, 113, 114, 114, 113, 117, 117, 104, 120, 121, 122, 122, 121, 125, 125, 120, 128, 128, 130, 130, 75, 133, 134, 135, 136, 136, 138, 138, 135, 141, 142, 142, 141, 145, 145, 134, 148, 149, 149, 151, 151, 148, 154, 155, 155, 154, 158, 158, 133, 161, 162, 163, 164, 164, 163, 162, 168, 169, 169, 168, 161, 173, 174, 175, 175, 174, 173, 179, 179, 0, 182, 183, 184, 185, 186, 187, 187, 189, 189, 186, 185, 193, 194, 194, 193, 197, 198, 198, 197, 201, 201, 184, 204, 205, 206, 206, 208, 208, 205, 211, 211, 213, 213, 204, 216, 217, 218, 218, 217, 216, 222, 222, 183, 225, 226, 226, 228, 229, 229, 231, 231, 228, 234, 235, 235, 234, 238, 238, 225, 241, 242, 243, 244, 244, 243, 247, 247, 242, 250, 251, 251, 250, 254, 254, 241, 257, 258, 259, 259, 258, 262, 262, 257, 265, 266, 266, 265, 269, 269, 182, 272, 273, 274, 275, 276, 276, 278, 278, 275, 274, 282, 282, 284, 285, 285, 284, 288, 288, 273, 291, 292, 293, 294, 294, 293, 297, 297, 292, 300, 301, 301, 300, 291, 305, 306, 306, 308, 308, 305, 311, 312, 312, 311, 272, 316, 317, 318, 318, 317, 321, 321, 323, 323, 325, 325, 316, 328, 329, 330, 331, 331, 330, 334, 334, 329, 337, 338, 338, 337, 341, 341, 328, 344, 345, 345, 347, 347, 344, 350, 351, 351, 350, 7, 7, 11, 11, 14, 14, 19, 19, 33, 33, 34, 34, 40, 40, 42, 42, 43, 43, 47, 47, 48, 48, 58, 58, 65, 65, 73, 73, 74, 74, 90, 90, 96, 96, 129, 129, 137, 137, 150, 150, 167, 167, 172, 172, 178, 178, 180, 180, 181, 181, 188, 188, 192, 192, 195, 195, 196, 196, 207, 207, 212, 212, 221, 221, 223, 223, 224, 224, 227, 227, 230, 230, 277, 277, 281, 281, 283, 283, 304, 304, 307, 307, 315, 315, 319, 319, 320, 320, 322, 322, 324, 324, 346, 346, 354, 354, 357, 357, 358, 358, 373, 373, 374, 374, 375, 375, 376, 376, 383, 383, 384, 384, 407, 407, 408, 408, 423, 423, 424, 424, 429, 429, 430, 430, 431, 431, 432, 432, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 463, 463, 464, 464, 465, 465, 466, 466, 471, 471, 472, 472, 473, 473, 474, 474),
                (-1, 0, 1, 2, 3, 4, 5, 6, 7, 7, 6, 10, 10, 5, 13, 14, 14, 13, 17, 17, 4, 20, 21, 22, 22, 21, 20, 26, 27, 27, 26, 30, 30, 3, 33, 33, 35, 35, 37, 38, 38, 37, 41, 41, 2, 44, 45, 46, 47, 47, 49, 49, 46, 52, 53, 53, 52, 56, 56, 45, 59, 60, 61, 61, 60, 59, 65, 65, 67, 67, 44, 70, 71, 71, 73, 73, 75, 75, 70, 78, 79, 79, 81, 81, 78, 84, 85, 85, 84, 88, 88, 1, 91, 92, 93, 94, 95, 96, 96, 95, 99, 99, 94, 102, 103, 103, 102, 106, 106, 93, 109, 110, 110, 109, 113, 113, 92, 116, 117, 117, 119, 120, 120, 119, 123, 123, 116, 126, 127, 128, 128, 127, 126, 132, 133, 133, 132, 91, 137, 138, 138, 140, 141, 142, 142, 141, 145, 145, 140, 148, 149, 149, 148, 137, 153, 154, 155, 156, 156, 155, 154, 160, 161, 161, 160, 153, 165, 166, 166, 168, 168, 165, 0, 172, 173, 174, 175, 176, 176, 178, 179, 179, 178, 182, 182, 175, 174, 186, 187, 188, 188, 190, 190, 187, 193, 193, 195, 195, 186, 198, 198, 200, 201, 201, 200, 204, 204, 173, 207, 208, 209, 210, 211, 211, 210, 209, 215, 216, 216, 215, 208, 220, 221, 221, 223, 223, 220, 226, 227, 227, 226, 230, 230, 207, 233, 234, 235, 235, 234, 238, 238, 240, 240, 233, 243, 243, 245, 245, 172, 248, 249, 249, 251, 252, 253, 254, 254, 253, 257, 257, 252, 260, 260, 251, 263, 264, 265, 265, 264, 268, 268, 263, 271, 271, 273, 273, 248, 276, 276, 278, 279, 280, 280, 282, 282, 279, 285, 286, 286, 285, 289, 289, 278, 292, 293, 294, 294, 293, 297, 297, 292, 300, 301, 301, 300, 25, 25, 34, 34, 36, 36, 48, 48, 64, 64, 66, 66, 72, 72, 74, 74, 80, 80, 111, 111, 112, 112, 114, 114, 115, 115, 118, 118, 131, 131, 136, 136, 139, 139, 152, 152, 159, 159, 164, 164, 167, 167, 171, 171, 177, 177, 185, 185, 189, 189, 194, 194, 199, 199, 214, 214, 219, 219, 222, 222, 236, 236, 237, 237, 239, 239, 244, 244, 246, 246, 247, 247, 250, 250, 261, 261, 262, 262, 272, 272, 277, 277, 281, 281, 304, 304, 307, 307, 308, 308, 309, 309, 310, 310, 317, 317, 318, 318, 331, 331, 332, 332, 337, 337, 338, 338, 347, 347, 348, 348, 349, 349, 350, 350, 351, 351, 352, 352, 357, 357, 358, 358, 371, 371, 372, 372, 377, 377, 378, 378, 385, 385, 386, 386, 391, 391, 392, 392, 393, 393, 394, 394, 407, 407, 408, 408, 409, 409, 410, 410, 419, 419, 420, 420, 421, 421, 422, 422, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 463, 463, 464, 464, 465, 465, 466, 466, 467, 467, 468, 468, 469, 469, 470, 470, 471, 471, 472, 472, 473, 473, 474, 474, 475, 475, 476, 476, 477, 477, 478, 478),
                (-1, 0, 1, 2, 3, 4, 5, 6, 6, 5, 4, 10, 11, 11, 10, 14, 15, 15, 14, 3, 19, 20, 20, 22, 23, 23, 22, 19, 27, 27, 29, 29, 31, 31, 2, 34, 35, 36, 37, 38, 38, 37, 41, 41, 36, 44, 45, 45, 44, 48, 48, 35, 51, 52, 53, 53, 52, 51, 57, 58, 58, 57, 34, 62, 63, 64, 64, 66, 66, 63, 69, 69, 71, 71, 62, 74, 75, 76, 76, 75, 79, 79, 74, 82, 82, 84, 84, 1, 87, 88, 89, 90, 91, 92, 92, 91, 90, 96, 97, 97, 96, 89, 101, 101, 103, 104, 104, 103, 107, 107, 88, 110, 111, 112, 113, 113, 112, 111, 117, 118, 118, 117, 121, 121, 110, 124, 125, 125, 127, 127, 124, 130, 131, 131, 130, 134, 134, 87, 137, 138, 139, 140, 140, 142, 142, 139, 138, 146, 146, 148, 149, 149, 148, 137, 153, 154, 155, 156, 156, 155, 159, 159, 154, 162, 162, 164, 164, 153, 167, 168, 169, 169, 168, 172, 172, 167, 0, 176, 177, 178, 179, 180, 181, 181, 183, 183, 180, 179, 187, 188, 188, 187, 191, 192, 192, 191, 195, 195, 178, 198, 199, 199, 201, 202, 202, 201, 205, 205, 198, 208, 209, 210, 210, 209, 213, 213, 208, 216, 216, 177, 219, 220, 221, 222, 223, 223, 222, 226, 226, 221, 229, 230, 230, 229, 233, 233, 220, 236, 237, 238, 238, 237, 236, 242, 243, 243, 242, 246, 246, 219, 249, 250, 251, 252, 252, 251, 255, 255, 250, 258, 259, 259, 258, 249, 263, 264, 265, 265, 264, 268, 268, 263, 271, 272, 272, 271, 275, 275, 176, 278, 279, 280, 281, 282, 283, 283, 282, 286, 286, 281, 289, 290, 290, 289, 293, 293, 280, 296, 297, 298, 298, 297, 296, 302, 303, 303, 302, 306, 306, 279, 309, 310, 310, 312, 312, 309, 315, 315, 317, 318, 318, 317, 321, 321, 278, 324, 324, 326, 327, 328, 329, 329, 328, 327, 333, 334, 334, 333, 326, 338, 339, 340, 340, 339, 343, 343, 338, 346, 346, 348, 348, 7, 7, 8, 8, 9, 9, 12, 12, 13, 13, 18, 18, 21, 21, 26, 26, 28, 28, 30, 30, 56, 56, 61, 61, 65, 65, 70, 70, 83, 83, 95, 95, 100, 100, 102, 102, 116, 116, 126, 126, 141, 141, 145, 145, 147, 147, 152, 152, 163, 163, 175, 175, 182, 182, 186, 186, 189, 189, 190, 190, 200, 200, 217, 217, 218, 218, 241, 241, 262, 262, 301, 301, 311, 311, 313, 313, 314, 314, 316, 316, 325, 325, 332, 332, 337, 337, 347, 347, 355, 355, 356, 356, 363, 363, 364, 364, 367, 367, 368, 368, 385, 385, 386, 386, 393, 393, 394, 394, 395, 395, 396, 396, 401, 401, 402, 402, 405, 405, 406, 406, 411, 411, 412, 412, 423, 423, 424, 424, 429, 429, 430, 430, 431, 431, 432, 432, 483, 483, 484, 484, 485, 485, 486, 486, 487, 487, 488, 488, 489, 489, 490, 490, 491, 491, 492, 492, 493, 493, 494, 494)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 2, 3, 4, 5, 6, 7, 7, 8, 8, 6, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 5, 6, 7, 8, 8, 7, 6, 7, 7, 3, 4, 5, 6, 6, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 8, 8, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 5, 2, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 8, 8, 3, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 5, 6, 7, 8, 8, 7, 6, 7, 7, 1, 2, 3, 4, 5, 6, 7, 7, 8, 8, 6, 5, 6, 7, 7, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 7, 3, 4, 5, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 2, 3, 4, 5, 6, 7, 7, 8, 8, 6, 5, 6, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 3, 4, 5, 6, 6, 5, 6, 6, 7, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8),
                (0, 1, 2, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 8, 8, 4, 5, 5, 6, 6, 7, 8, 8, 7, 8, 8, 3, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 7, 8, 8, 4, 5, 6, 6, 7, 7, 8, 8, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 2, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 7, 6, 7, 7, 4, 5, 6, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 3, 4, 5, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 5, 6, 7, 7, 8, 8, 6, 1, 2, 3, 4, 5, 6, 6, 7, 8, 8, 7, 8, 8, 5, 4, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 8, 5, 6, 6, 7, 8, 8, 7, 8, 8, 3, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 7, 6, 7, 7, 8, 8, 5, 6, 6, 7, 7, 2, 3, 4, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 8, 8, 3, 4, 4, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 6, 6, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 5, 5, 8, 8, 8, 8, 8, 8, 5, 5, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 6, 6, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8),
                (0, 1, 2, 3, 4, 5, 6, 7, 7, 6, 5, 6, 7, 7, 6, 7, 8, 8, 7, 4, 5, 6, 6, 7, 8, 8, 7, 5, 6, 6, 7, 7, 8, 8, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 4, 5, 6, 7, 7, 8, 8, 6, 7, 7, 8, 8, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 8, 8, 2, 3, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 5, 6, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 3, 4, 5, 6, 7, 7, 8, 8, 6, 5, 6, 6, 7, 8, 8, 7, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 8, 8, 5, 6, 7, 8, 8, 7, 8, 8, 6, 1, 2, 3, 4, 5, 6, 7, 7, 8, 8, 6, 5, 6, 7, 7, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 2, 3, 4, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 8, 8, 7, 8, 8, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 8, 8, 4, 5, 6, 6, 7, 7, 5, 6, 6, 7, 8, 8, 7, 8, 8, 3, 4, 4, 5, 6, 7, 8, 8, 7, 6, 7, 8, 8, 7, 5, 6, 7, 8, 8, 7, 8, 8, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 5, 5, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((9, 10, 16, 17, 21, 22, 27, 28, 30, 31, 38, 39, 52, 53, 55, 56, 60, 61, 67, 68, 71, 72, 81, 82, 84, 85, 88, 89, 94, 95, 99, 100, 102, 103, 108, 109, 111, 112, 115, 116, 118, 119, 123, 124, 126, 127, 131, 132, 139, 140, 143, 144, 146, 147, 152, 153, 156, 157, 159, 160, 165, 166, 170, 171, 176, 177, 190, 191, 199, 200, 202, 203, 209, 210, 214, 215, 219, 220, 232, 233, 236, 237, 239, 240, 245, 246, 248, 249, 252, 253, 255, 256, 260, 261, 263, 264, 267, 268, 270, 271, 279, 280, 286, 287, 289, 290, 295, 296, 298, 299, 302, 303, 309, 310, 313, 314, 326, 327, 332, 333, 335, 336, 339, 340, 342, 343, 348, 349, 352, 353, 355, 356, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 377, 378, 379, 380, 381, 382, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 425, 426, 427, 428, 433, 434, 435, 436, 437, 438, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 467, 468, 469, 470, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510),
                (8, 9, 11, 12, 15, 16, 18, 19, 23, 24, 28, 29, 31, 32, 39, 40, 42, 43, 50, 51, 54, 55, 57, 58, 62, 63, 68, 69, 76, 77, 82, 83, 86, 87, 89, 90, 97, 98, 100, 101, 104, 105, 107, 108, 121, 122, 124, 125, 129, 130, 134, 135, 143, 144, 146, 147, 150, 151, 157, 158, 162, 163, 169, 170, 180, 181, 183, 184, 191, 192, 196, 197, 202, 203, 205, 206, 212, 213, 217, 218, 224, 225, 228, 229, 231, 232, 241, 242, 255, 256, 258, 259, 266, 267, 269, 270, 274, 275, 283, 284, 287, 288, 290, 291, 295, 296, 298, 299, 302, 303, 305, 306, 311, 312, 313, 314, 315, 316, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 333, 334, 335, 336, 339, 340, 341, 342, 343, 344, 345, 346, 353, 354, 355, 356, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 373, 374, 375, 376, 379, 380, 381, 382, 383, 384, 387, 388, 389, 390, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 411, 412, 413, 414, 415, 416, 417, 418, 423, 424, 425, 426, 427, 428, 429, 430, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510),
                (16, 17, 24, 25, 32, 33, 39, 40, 42, 43, 46, 47, 49, 50, 54, 55, 59, 60, 67, 68, 72, 73, 77, 78, 80, 81, 85, 86, 93, 94, 98, 99, 105, 106, 108, 109, 114, 115, 119, 120, 122, 123, 128, 129, 132, 133, 135, 136, 143, 144, 150, 151, 157, 158, 160, 161, 165, 166, 170, 171, 173, 174, 184, 185, 193, 194, 196, 197, 203, 204, 206, 207, 211, 212, 214, 215, 224, 225, 227, 228, 231, 232, 234, 235, 239, 240, 244, 245, 247, 248, 253, 254, 256, 257, 260, 261, 266, 267, 269, 270, 273, 274, 276, 277, 284, 285, 287, 288, 291, 292, 294, 295, 299, 300, 304, 305, 307, 308, 319, 320, 322, 323, 330, 331, 335, 336, 341, 342, 344, 345, 349, 350, 351, 352, 353, 354, 357, 358, 359, 360, 361, 362, 365, 366, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 387, 388, 389, 390, 391, 392, 397, 398, 399, 400, 403, 404, 407, 408, 409, 410, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 425, 426, 427, 428, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, -2, 1, 1, 1, 1, 0, 0, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, -2, 0, -2, -2, 1, 1, 1, 2, 0, 2, -2, 2, -2, 2, 2, -2, 0, 0, 1, -2, 2, 0, -2, -2, 1, 2, -2, 2, 0, 0, -2, -2, -2, -2, 0, 0, 0, -2, 0, -2, 0, -2, -2, -2, 0, 0, -2, 1, -2, -2, -2, 1, 1, -2, -2, 2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, 1, 0, -2, -2, -2, 2, -2, -2, -2, 0, -2, -2, -2, -2, 2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, 1, 1, 0, -2, -2, -2, -2, 0, -2, -2, 2, 1, -2, -2, -2, -2, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, 2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 0, 2, 0, -2, 0, 0, 1, 1, 1, 2, 1, 1, -2, 2, 0, 0, 2, 0, 1, 1, 2, 0, 0, 0, 1, 0, 1, 2, 1, 2, 0, 1, 1, 0, 1, 1, 0, 0, -2, -2, 1, 1, -2, -2, 1, 1, 2, 1, 0, -2, 0, 2, 2, 1, 1, -2, 0, -2, 1, -2, -2, -2, -2, -2, -2, -2, 1, 0, -2, -2, 0, 0, 1, 2, -2, 2, -2, -2, -2, -2, 1, 2, 0, -2, -2, -2, 1, 0, 1, 1, -2, -2, 2, 1, -2, -2, -2, 1, -2, -2, 0, 0, 0, 0, 2, 2, -2, -2, 0, -2, -2, -2, -2, -2, 1, 1, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, 0, -2, -2, -2, -2, 2, -2, -2, -2, -2, 0, 0, -2, -2, -2, -2, 1, 0, -2, 2, 0, -2, 1, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 0, 0, 1, 2, -2, -2, 1, -2, -2, -2, 1, 0, -2, -2, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, 1, -2, -2, -2, -2, -2, 1, 1, -2, -2, -2, -2, -2, -2, 0, 0, -2, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, 0, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, 1, -2, -2, 2, -2, -2, 1, -2, -2, 2, 0, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 1, 1, -2, -2, 0, 0, 0, 1, 1, 2, 1, 1, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, 0, 1, 2, 1, 0, -2, 2, 0, -2, -2, -2, -2, -2, 1, 0, 1, 2, -2, -2, 0, 1, -2, -2, -2, -2, 2, 2, -2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((29516454, 968977, 44568188, 8413001, 15744038, 540558, 795582, 11881806, 1371414, 1525456, 45940494, 1416839, 56033, 56033, 68567, 3152512, 5031608, 258141, 405509, 36800210, 34146544, 9078326, 13746256, 1591456, 24316919, 68567, -131072, 1108281, 1251232, 1535980, 1656718, 22087124, 19096339, 68567, 1357138, 1154520, 1256733, 641936, 724037, 1077416, 1141954, 757667, 1912893, 103290, 195145, 68567, 83804, 1641747, 46858, 18649150, 18464894, 24185218, 28230463, 1404997, 56033, 18410685, 20310496, 1205042, 1321827, -131072, 4585107, -131072, -131072, 1691649, 1737312, 493669, 46858, 23214072, 46858, -131072, 68567, -131072, 46858, 68567, -131072, 11293262, 9325304, 1651450, -131072, 46858, 33304979, -131072, -131072, 906697, 46858, -131072, 83804, 6556334, 6054382, -131072, -131072, -131072, -131072, 41277348, 41966276, 13754473, -131072, 32805027, -131072, 31741048, -131072, -131072, -131072, 34169206, 32181741, -131072, 1776994, -131072, -131072, -131072, 407537, 1810316, -131072, -131072, 46858, -131072, -131072, -131072, -131072, -131072, -131072, 8405652, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 800229, 7188240, -131072, -131072, -131072, 68567, -131072, -131072, -131072, 39660190, -131072, -131072, -131072, -131072, 83804, -131072, -131072, 14708472, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1003515, 1108356, 13116422, -131072, -131072, -131072, -131072, 3793179, -131072, -131072, 83804, 953245, -131072, -131072, -131072, -131072, 56033, 712572, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 46858, -131072, 56033, -131072, -131072, -131072, -131072, -131072, 20509651, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 32236968, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072),
                (27391894, 724503, 37406376, 5284170, 17720116, 212233, 7247426, 1513009, 44566694, 1377766, 68567, 954422, 1257289, 1160222, 83804, 56033, 28448155, 983040, 3904877, 542684, 1273713, 1442091, 1597524, 19090289, 23497959, 9834861, 13695944, 7870195, 46858, 596689, 7975306, 529280, 68567, 19017009, 56033, 23021487, -131072, 13700419, 11796034, 352183, 488099, 447821, 68567, 764145, 924930, -131072, 46858, 31464166, 28091446, 46858, 24002226, 1679350, 1799131, 68567, 26204547, 25456269, 18939147, 1706121, 45999286, 1630766, 46858, 1711320, 56033, 30693485, 1465182, 1587548, 33489500, 1647137, 1897566, 27613098, 32202178, -131072, -131072, 871412, 944910, -131072, -131072, 1076796, 1174373, 68567, 1351620, 17159495, -131072, 7097632, 68567, 56033, 827260, 1468840, -131072, 39417192, -131072, 1805922, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 643538, 5801802, -131072, -131072, 34060482, 33391925, 1516343, 46858, -131072, 46858, -131072, -131072, -131072, -131072, 1569725, 46858, 42621406, -131072, -131072, -131072, 584895, 5565259, 531717, 559585, -131072, -131072, 83804, 1398125, -131072, -131072, -131072, 110463, -131072, -131072, 2237185, 3113596, 1952471, 2737676, 68567, 68567, -131072, -131072, 38658984, -131072, -131072, -131072, -131072, -131072, 1097308, 1139890, 1064529, 46858, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1844363, -131072, 28255106, -131072, -131072, -131072, -131072, 46858, -131072, -131072, -131072, -131072, 32108153, 34050064, -131072, -131072, -131072, -131072, 620428, 8648233, -131072, 56033, 7312861, -131072, 1855224, -131072, -131072, -131072, 27483458, -131072, -131072, -131072, -131072, -131072, 1398461, 30808174, -131072, -131072, -131072, -131072, -131072, -131072, 6698962, -131072, -131072, -131072, 9965244, 11789584, 960514, 68567, -131072, -131072, 164097, -131072, -131072, -131072, 1709805, 40583236, -131072, -131072, 1603726, 46858, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 28018870, -131072, 1505389, -131072, -131072, -131072, -131072, -131072, 393178, 440117, -131072, -131072, -131072, -131072, -131072, -131072, 6553306, 7106472, -131072, -131072, -131072, -131072, -131072, 40610238, -131072, -131072, -131072, 1571247, -131072, 38985640, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 11791142, -131072, -131072, 667848, -131072, -131072, 67011, -131072, -131072, 1770367, -131072, -131072, 46858, 44927686, -131072, -131072, -131072, -131072, -131072, -131072, 1140098, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072),
                (30235935, 759528, 38658048, 7119044, 20914772, 254422, 7958326, 1538414, 44577396, 1430581, 56033, 1079846, 1324561, 1252578, 68567, 1647216, 68567, 1359537, 3804826, 750555, 1632322, 1461441, 1609813, -131072, -131072, 13200494, 18287654, 9688893, 985525, 1196157, 56033, 325724, 477841, -131072, -131072, -131072, -131072, -131072, -131072, 33068504, -131072, -131072, -131072, -131072, -131072, 1696361, 46055012, 1599630, 46858, 1751147, 39380402, -131072, 46858, 33434543, -131072, -131072, -131072, -131072, -131072, 646170, 8645402, 632178, 56033, -131072, -131072, 14467401, 1237636, -131072, -131072, -131072, -131072, 46858, 46858, -131072, -131072, -131072, 46858, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 713639, 757558, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1748918, -131072, -131072, 46858, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((17447, 8188, 21568, 15251, 3208, 6691, 21090, 424, 7781, 20028, 21842, 21776, 13223, 16132, 3493, 12688, 1633, 4737, 20450, 7005, 20489, 21830, 17916, 1167, 8397, 9570, 21845, 38, 1834, 4515, 18341, 11479, 20127, 6629, 134, 5980, 18423, 131, 4427, 2101, 18116, 10353, 1079, 1755, 20080, 10992, 898, 2828, 12927, 14487, 1464, 2604, 82, 385, 6860, 12136, 2052, 16447, 21736, 21845, 17006, 2893, 17554, 7459, 20006, 7982, 21433, 21538, 12525, 21845, 11852, 21845, 20837, 17847, 21845, 6320, 19704, 11818, 21845, 7986, 607, 2849, 18153, 1748, 14070, 21845, 13949, 6399, 18832, 3197, 18548, 203, 4755, 16257, 2731, 5601, 0, 16991, 21845, 4369, 21845, 5174, 20074, 2683, 16384, 21845, 6162, 1481, 13653, 0, 3149, 21631, 21845, 21845, 12136, 7437, 0, 533, 11218, 9362, 19946, 252, 0, 21845, 14564, 12578, 0, 10082, 20436, 271, 3932, 4915, 0, 0, 927, 5749, 18022, 21845, 16705, 8402, 21845, 2149, 65, 759, 0, 0, 5749, 11398, 21845, 10280, 21845, 0, 2849, 0, 2832, 21337, 14564, 5041, 19325, 1150, 12743, 563, 0, 0, 2664, 14043, 21845, 15124, 21845, 0, 819, 21370, 21845, 520, 8738, 0, 21845, 11498, 1092, 643, 12483, 19661, 0, 809, 6722, 0, 1351, 21845, 16991, 3013, 0, 0, 2789, 21845, 21092, 19859, 21845, 0, 2731, 923, 0, 17476, 21845, 19418, 21845, 9709, 1456, 2913, 16384, 0, 8192, 10923, 21845, 21845, 19859, 5461, 10923, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 0, 0, 21845, 21845, 0, 0, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 10923, 10923, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845),
                (14203, 4389, 21025, 13546, 1942, 3314, 20925, 15980, 21713, 21279, 5421, 796, 5896, 19405, 2138, 2121, 21148, 11265, 1654, 1893, 21526, 1332, 8912, 19546, 3361, 3473, 334, 604, 15869, 14731, 21717, 20590, 3013, 21286, 13623, 6756, 21845, 8162, 18958, 670, 6497, 20285, 2110, 2466, 20339, 21845, 16432, 7282, 21544, 2874, 20805, 1142, 15066, 4031, 587, 2570, 18933, 20202, 21840, 21590, 10194, 1365, 18946, 2427, 16991, 1118, 6314, 3099, 20480, 16880, 551, 1564, 10114, 14303, 21693, 21255, 8831, 97, 1332, 7443, 500, 3351, 21845, 110, 3841, 624, 14564, 9709, 21845, 13222, 21845, 3641, 21845, 2226, 12647, 19418, 0, 21845, 9102, 1181, 13443, 0, 21845, 4450, 533, 1066, 15124, 21845, 14312, 19661, 4855, 8738, 21845, 21803, 17828, 5958, 21845, 17476, 1150, 4855, 18569, 364, 5851, 19661, 2849, 2120, 83, 910, 15604, 0, 5680, 21845, 0, 2630, 212, 686, 17476, 336, 2608, 1285, 9866, 3449, 21845, 10194, 21845, 5461, 21845, 18504, 21798, 21504, 9362, 0, 19661, 0, 21845, 824, 7598, 10923, 21845, 125, 6827, 16147, 21845, 18569, 0, 5461, 19418, 21845, 13107, 0, 21845, 13107, 0, 20480, 11916, 4369, 18204, 3799, 0, 19357, 21812, 21845, 9557, 3972, 21845, 21141, 0, 21845, 10923, 19546, 0, 21845, 2185, 117, 1248, 1425, 8192, 21845, 3641, 0, 5041, 7282, 575, 3799, 0, 2081, 21845, 540, 32, 26, 2819, 143, 15226, 16384, 21845, 21845, 0, 7282, 1030, 0, 21845, 107, 1365, 158, 3745, 6242, 560, 10923, 20560, 0, 5958, 21845, 14564, 0, 2131, 14564, 21845, 18725, 21845, 20165, 0, 21845, 10923, 16384, 21845, 58, 879, 8738, 400, 918, 0, 2427, 0, 20, 950, 21845, 767, 21845, 17476, 0, 1791, 21845, 1456, 21845, 20805, 0, 21141, 17873, 21845, 21845, 18725, 1456, 0, 0, 261, 21845, 235, 21083, 21845, 21845, 8738, 0, 21845, 21566, 21845, 21845, 14043, 3641, 21845, 21845, 0, 560, 0, 21845, 21005, 0, 21845, 520, 0, 0, 428, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845),
                (12030, 3568, 21050, 11437, 1651, 3070, 21472, 15296, 21705, 21380, 5334, 759, 6086, 19727, 2305, 1216, 16549, 10037, 1584, 1932, 21489, 803, 8584, 18380, 4356, 2590, 272, 882, 17005, 21276, 11967, 376, 4791, 21354, 1726, 166, 4645, 20537, 11327, 10824, 21845, 6899, 21845, 4073, 18485, 19868, 21837, 21636, 9264, 984, 20753, 21845, 16384, 6604, 21845, 3576, 248, 1409, 20025, 16434, 21747, 21565, 3523, 588, 10037, 124, 1630, 9261, 1015, 0, 18204, 3722, 531, 1126, 10348, 21845, 17970, 9198, 21845, 21716, 18046, 12483, 21845, 2087, 177, 30, 580, 15604, 21845, 19806, 21823, 21845, 4855, 0, 1266, 3013, 266, 21845, 16384, 21435, 21845, 21845, 16182, 2731, 21845, 21834, 20025, 18380, 18380, 4356, 4356, 21354, 21354, 1726, 1726, 166, 166, 4645, 4645, 20537, 20537, 11327, 11327, 21845, 21845, 6899, 6899, 21845, 21845, 4073, 4073, 18485, 18485, 21845, 21845, 21845, 21845, 3576, 3576, 248, 248, 1409, 1409, 20025, 20025, 588, 588, 10037, 10037, 9261, 9261, 1015, 1015, 0, 0, 18204, 18204, 1126, 1126, 10348, 10348, 21845, 21845, 9198, 9198, 21845, 21845, 21716, 21716, 18046, 18046, 12483, 12483, 21845, 21845, 2087, 2087, 177, 177, 30, 30, 580, 580, 15604, 15604, 21845, 21845, 21845, 21845, 4855, 4855, 0, 0, 1266, 1266, 3013, 3013, 266, 266, 21845, 21845, 16384, 16384, 21845, 21845, 21845, 21845, 2731, 2731, 21845, 21845, 21834, 21834, 20025, 20025, 18380, 18380, 18380, 18380, 4356, 4356, 4356, 4356, 21354, 21354, 21354, 21354, 1726, 1726, 1726, 1726, 166, 166, 166, 166, 4645, 4645, 4645, 4645, 20537, 20537, 20537, 20537, 11327, 11327, 11327, 11327, 21845, 21845, 21845, 21845, 6899, 6899, 6899, 6899, 21845, 21845, 21845, 21845, 4073, 4073, 4073, 4073, 18485, 18485, 18485, 18485, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 3576, 3576, 3576, 3576, 248, 248, 248, 248, 1409, 1409, 1409, 1409, 20025, 20025, 20025, 20025, 588, 588, 588, 588, 10037, 10037, 10037, 10037, 9261, 9261, 9261, 9261, 1015, 1015, 1015, 1015, 0, 0, 0, 0, 18204, 18204, 18204, 18204, 1126, 1126, 1126, 1126, 10348, 10348, 10348, 10348, 21845, 21845, 21845, 21845, 9198, 9198, 9198, 9198, 21845, 21845, 21845, 21845, 21716, 21716, 21716, 21716, 18046, 18046, 18046, 18046, 12483, 12483, 12483, 12483, 21845, 21845, 21845, 21845, 2087, 2087, 2087, 2087, 177, 177, 177, 177, 30, 30, 30, 30, 580, 580, 580, 580, 15604, 15604, 15604, 15604, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 4855, 4855, 4855, 4855, 0, 0, 0, 0, 1266, 1266, 1266, 1266, 3013, 3013, 3013, 3013, 266, 266, 266, 266, 21845, 21845, 21845, 21845, 16384, 16384, 16384, 16384, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 2731, 2731, 2731, 2731, 21845, 21845, 21845, 21845, 21834, 21834, 21834, 21834, 20025, 20025, 20025, 20025, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 9, 5, 7, 15, 21, 27, 13, 11, 111, 71, 19, 31, 23, 17, 37, 41, 59, 47, 73, 171, 25, 51, 29, 75, 217, 121, 33, 55, 85, 35, 57, 39, 143, 49, 67, 161, 45, 95, 155, 43, 109, 131, 123, 87, 129, 79, 63, 119, 151, 53, 169, 141, 61, 81, 91, 69, 193, 219, 65, -1, -1, 93, 137, 125, 203, 195, 101, 221, 89, 223, 97, 77, 225, 83, 165, 105, 227, 103, 185, -1, -1, 189, 135, 229, 127, 107, 167, -1, -1, -1, -1, 147, 183, 117, 231, 99, 233, 209, 235, -1, -1, 173, 149, 237, 177, -1, -1, 239, 115, 113, 241, 243, 175, -1, -1, -1, -1, -1, -1, 133, 245, -1, -1, -1, -1, -1, -1, 199, 159, -1, -1, 247, 153, -1, -1, 249, 139, -1, -1, -1, -1, 145, 251, 253, 207, -1, -1, -1, -1, -1, -1, 255, 205, 213, 157, -1, -1, -1, -1, 163, 257, 259, 179, 181, 261, -1, -1, 263, 197, 187, 265, -1, -1, 267, 269, -1, -1, -1, -1, -1, -1, -1, -1, 271, 191, 273, 211, -1, -1, -1, -1, 275, 201, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 277, 215, 279, 281, -1, -1, -1, -1, 283, 285, 287, 289, -1, -1, 291, 293, 295, 297, 299, 301, -1, -1, -1, -1, 303, 305, 307, 309, -1, -1, -1, -1, 311, 313, 315, 317, 319, 321, 323, 325, -1, -1, 327, 329, -1, -1, -1, -1, 331, 333, -1, -1, -1, -1, -1, -1, 335, 337, 339, 341, 343, 345, -1, -1, 347, 349, -1, -1, -1, -1, -1, -1, -1, -1, 351, 353, 355, 357, -1, -1, -1, -1, 359, 361, 363, 365, 367, 369, 371, 373, -1, -1, -1, -1, 375, 377, 379, 381, -1, -1, -1, -1, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 407, 409, 411, 413, 415, 417, 419, 421, 423, 425, 427, 429, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 431, 433, 435, 437, 439, 441, 443, 445, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 447, 449, 451, 453, 455, 457, 459, 461, 463, 465, 467, 469, 471, 473, 475, 477, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 11, 17, 29, 9, 57, 45, 15, 25, 13, 33, 21, 65, 161, 19, 39, 129, 213, 53, 23, 87, 51, 27, 77, 83, 37, 31, 179, 107, 99, 147, 35, 49, 301, 43, 73, 133, 41, 167, 121, 117, 187, 303, 47, 63, 237, 155, 243, 177, 109, 55, 137, 71, 111, 59, 283, 113, 61, 217, 89, 195, 173, 103, 67, 69, 185, 165, 199, -1, -1, 75, 269, -1, -1, 207, 79, 81, 125, 93, 305, 253, 85, 233, 97, 95, 307, 91, 309, 171, 311, -1, -1, -1, -1, -1, -1, 203, 101, 313, 315, 105, 221, 201, 143, 317, 119, -1, -1, -1, -1, 263, 115, 141, 319, -1, -1, 153, 145, 251, 123, -1, -1, 127, 249, -1, -1, 321, 131, 323, 325, 135, 245, 159, 157, 193, 139, -1, -1, 229, 327, -1, -1, -1, -1, 149, 293, 257, 151, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 163, 329, 189, 331, -1, -1, 333, 169, -1, -1, -1, -1, 235, 175, -1, -1, -1, -1, 181, 277, 335, 183, 191, 337, 231, 339, -1, -1, 227, 341, -1, -1, -1, -1, 225, 197, -1, -1, -1, -1, -1, -1, 205, 343, -1, -1, 209, 273, 297, 211, -1, -1, 215, 345, 347, 349, 219, 259, 351, 353, 271, 223, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 239, 355, 241, 357, -1, -1, -1, -1, 291, 247, -1, -1, -1, -1, -1, -1, 299, 255, -1, -1, -1, -1, 359, 261, -1, -1, 361, 265, 363, 267, -1, -1, -1, -1, -1, -1, 365, 275, -1, -1, 279, 367, 369, 281, -1, -1, 285, 371, 373, 287, 289, 375, 377, 379, -1, -1, 381, 295, -1, -1, -1, -1, -1, -1, 383, 385, 387, 389, -1, -1, -1, -1, 391, 393, -1, -1, -1, -1, -1, -1, 395, 397, 399, 401, 403, 405, -1, -1, -1, -1, -1, -1, 407, 409, 411, 413, -1, -1, 415, 417, -1, -1, -1, -1, -1, -1, -1, -1, 419, 421, -1, -1, -1, -1, -1, -1, -1, -1, 423, 425, -1, -1, -1, -1, 427, 429, -1, -1, -1, -1, 431, 433, -1, -1, 435, 437, 439, 441, 443, 445, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 447, 449, 451, 453, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 455, 457, 459, 461, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 463, 465, 467, 469, 471, 473, 475, 477, -1, -1, -1, -1, 479, 481, 483, 485, 487, 489, 491, 493, -1, -1, -1, -1, -1, -1, -1, -1, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 11, 17, 59, 9, 45, 51, 15, 25, 13, 29, 21, 71, 39, 19, 31, 63, 81, 55, 23, 107, 109, 27, 65, 35, 37, 79, 41, 83, 33, 111, 113, 115, 117, 119, 121, 43, 123, 125, 127, 129, 131, 47, 99, 75, 49, 95, 87, 133, 53, 57, 135, 137, 139, 141, 143, 61, 89, 97, 69, 145, 147, 85, 67, 149, 151, 153, 155, 73, 93, 157, 159, 161, 77, 163, 165, 167, 169, 171, 173, 175, 177, 179, 181, 183, 185, 91, 105, 187, 189, 191, 193, 195, 197, 199, 201, 101, 203, 205, 103, 207, 209, 211, 213, 215, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 237, 239, 241, 243, 245, 247, 249, 251, 253, 255, 257, 259, 261, 263, 265, 267, 269, 271, 273, 275, 277, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 341, 343, 345, 347, 349, 351, 353, 355, 357, 359, 361, 363, 365, 367, 369, 371, 373, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 415, 417, 419, 421, 423, 425, 427, 429, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 431, 433, 435, 437, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 439, 441, 443, 445, 447, 449, 451, 453, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 455, 457, 459, 461, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 463, 465, 467, 469, 471, 473, 475, 477, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 479, 481, 483, 485, 487, 489, 491, 493, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 495, 497, 499, 501, 503, 505, 507, 509, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 10, 6, 8, 16, 22, 28, 14, 12, 112, 72, 20, 32, 24, 18, 38, 42, 60, 48, 74, 172, 26, 52, 30, 76, 218, 122, 34, 56, 86, 36, 58, 40, 144, 50, 68, 162, 46, 96, 156, 44, 110, 132, 124, 88, 130, 80, 64, 120, 152, 54, 170, 142, 62, 82, 92, 70, 194, 220, 66, -1, -1, 94, 138, 126, 204, 196, 102, 222, 90, 224, 98, 78, 226, 84, 166, 106, 228, 104, 186, -1, -1, 190, 136, 230, 128, 108, 168, -1, -1, -1, -1, 148, 184, 118, 232, 100, 234, 210, 236, -1, -1, 174, 150, 238, 178, -1, -1, 240, 116, 114, 242, 244, 176, -1, -1, -1, -1, -1, -1, 134, 246, -1, -1, -1, -1, -1, -1, 200, 160, -1, -1, 248, 154, -1, -1, 250, 140, -1, -1, -1, -1, 146, 252, 254, 208, -1, -1, -1, -1, -1, -1, 256, 206, 214, 158, -1, -1, -1, -1, 164, 258, 260, 180, 182, 262, -1, -1, 264, 198, 188, 266, -1, -1, 268, 270, -1, -1, -1, -1, -1, -1, -1, -1, 272, 192, 274, 212, -1, -1, -1, -1, 276, 202, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 278, 216, 280, 282, -1, -1, -1, -1, 284, 286, 288, 290, -1, -1, 292, 294, 296, 298, 300, 302, -1, -1, -1, -1, 304, 306, 308, 310, -1, -1, -1, -1, 312, 314, 316, 318, 320, 322, 324, 326, -1, -1, 328, 330, -1, -1, -1, -1, 332, 334, -1, -1, -1, -1, -1, -1, 336, 338, 340, 342, 344, 346, -1, -1, 348, 350, -1, -1, -1, -1, -1, -1, -1, -1, 352, 354, 356, 358, -1, -1, -1, -1, 360, 362, 364, 366, 368, 370, 372, 374, -1, -1, -1, -1, 376, 378, 380, 382, -1, -1, -1, -1, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 432, 434, 436, 438, 440, 442, 444, 446, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 12, 18, 30, 10, 58, 46, 16, 26, 14, 34, 22, 66, 162, 20, 40, 130, 214, 54, 24, 88, 52, 28, 78, 84, 38, 32, 180, 108, 100, 148, 36, 50, 302, 44, 74, 134, 42, 168, 122, 118, 188, 304, 48, 64, 238, 156, 244, 178, 110, 56, 138, 72, 112, 60, 284, 114, 62, 218, 90, 196, 174, 104, 68, 70, 186, 166, 200, -1, -1, 76, 270, -1, -1, 208, 80, 82, 126, 94, 306, 254, 86, 234, 98, 96, 308, 92, 310, 172, 312, -1, -1, -1, -1, -1, -1, 204, 102, 314, 316, 106, 222, 202, 144, 318, 120, -1, -1, -1, -1, 264, 116, 142, 320, -1, -1, 154, 146, 252, 124, -1, -1, 128, 250, -1, -1, 322, 132, 324, 326, 136, 246, 160, 158, 194, 140, -1, -1, 230, 328, -1, -1, -1, -1, 150, 294, 258, 152, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 164, 330, 190, 332, -1, -1, 334, 170, -1, -1, -1, -1, 236, 176, -1, -1, -1, -1, 182, 278, 336, 184, 192, 338, 232, 340, -1, -1, 228, 342, -1, -1, -1, -1, 226, 198, -1, -1, -1, -1, -1, -1, 206, 344, -1, -1, 210, 274, 298, 212, -1, -1, 216, 346, 348, 350, 220, 260, 352, 354, 272, 224, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 240, 356, 242, 358, -1, -1, -1, -1, 292, 248, -1, -1, -1, -1, -1, -1, 300, 256, -1, -1, -1, -1, 360, 262, -1, -1, 362, 266, 364, 268, -1, -1, -1, -1, -1, -1, 366, 276, -1, -1, 280, 368, 370, 282, -1, -1, 286, 372, 374, 288, 290, 376, 378, 380, -1, -1, 382, 296, -1, -1, -1, -1, -1, -1, 384, 386, 388, 390, -1, -1, -1, -1, 392, 394, -1, -1, -1, -1, -1, -1, 396, 398, 400, 402, 404, 406, -1, -1, -1, -1, -1, -1, 408, 410, 412, 414, -1, -1, 416, 418, -1, -1, -1, -1, -1, -1, -1, -1, 420, 422, -1, -1, -1, -1, -1, -1, -1, -1, 424, 426, -1, -1, -1, -1, 428, 430, -1, -1, -1, -1, 432, 434, -1, -1, 436, 438, 440, 442, 444, 446, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 448, 450, 452, 454, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 456, 458, 460, 462, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 464, 466, 468, 470, 472, 474, 476, 478, -1, -1, -1, -1, 480, 482, 484, 486, 488, 490, 492, 494, -1, -1, -1, -1, -1, -1, -1, -1, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 12, 18, 60, 10, 46, 52, 16, 26, 14, 30, 22, 72, 40, 20, 32, 64, 82, 56, 24, 108, 110, 28, 66, 36, 38, 80, 42, 84, 34, 112, 114, 116, 118, 120, 122, 44, 124, 126, 128, 130, 132, 48, 100, 76, 50, 96, 88, 134, 54, 58, 136, 138, 140, 142, 144, 62, 90, 98, 70, 146, 148, 86, 68, 150, 152, 154, 156, 74, 94, 158, 160, 162, 78, 164, 166, 168, 170, 172, 174, 176, 178, 180, 182, 184, 186, 92, 106, 188, 190, 192, 194, 196, 198, 200, 202, 102, 204, 206, 104, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 432, 434, 436, 438, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 440, 442, 444, 446, 448, 450, 452, 454, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 456, 458, 460, 462, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 464, 466, 468, 470, 472, 474, 476, 478, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 480, 482, 484, 486, 488, 490, 492, 494, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 496, 498, 500, 502, 504, 506, 508, 510, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 8, 8, 5, 5, 15, 15, 12, 12, 6, 6, 14, 14, 22, 22, 7, 7, 24, 24, 13, 13, 28, 28, 31, 31, 16, 16, 33, 33, 17, 17, 41, 41, 38, 38, 19, 19, 35, 35, 23, 23, 51, 51, 29, 29, 32, 32, 18, 18, 54, 54, 48, 48, 60, 60, 36, 36, 57, 57, 11, 11, 20, 20, 25, 25, 73, 73, 47, 47, 55, 55, 75, 75, 30, 30, 45, 45, 70, 70, 56, 56, 63, 63, 39, 39, 72, 72, 97, 97, 68, 68, 79, 79, 77, 77, 87, 87, 42, 42, 10, 10, 111, 111, 110, 110, 95, 95, 49, 49, 27, 27, 44, 44, 65, 65, 86, 86, 46, 46, 43, 43, 121, 121, 84, 84, 64, 64, 138, 138, 53, 53, 34, 34, 143, 143, 93, 93, 104, 104, 50, 50, 134, 134, 40, 40, 156, 156, 130, 130, 37, 37, 161, 161, 76, 76, 88, 88, 52, 52, 21, 21, 103, 103, 114, 114, 106, 106, 164, 164, 165, 165, 94, 94, 80, 80, 171, 171, 83, 83, 186, 186, 58, 58, 67, 67, 170, 170, 129, 129, 194, 194, 66, 66, 154, 154, 146, 146, 99, 99, 188, 188, 155, 155, 210, 210, 26, 26, 59, 59, 69, 69, 71, 71, 74, 74, 78, 78, 85, 85, 96, 96, 98, 98, 100, 100, 105, 105, 109, 109, 112, 112, 113, 113, 122, 122, 133, 133, 137, 137, 144, 144, 145, 145, 153, 153, 162, 162, 163, 163, 166, 166, 169, 169, 172, 172, 175, 175, 176, 176, 185, 185, 187, 187, 193, 193, 209, 209, 211, 211, 212, 212, 217, 217, 218, 218, 219, 219, 220, 220, 223, 223, 224, 224, 225, 225, 226, 226, 227, 227, 228, 228, 233, 233, 234, 234, 235, 235, 236, 236, 241, 241, 242, 242, 243, 243, 244, 244, 245, 245, 246, 246, 247, 247, 248, 248, 251, 251, 252, 252, 257, 257, 258, 258, 265, 265, 266, 266, 267, 267, 268, 268, 269, 269, 270, 270, 273, 273, 274, 274, 283, 283, 284, 284, 285, 285, 286, 286, 291, 291, 292, 292, 293, 293, 294, 294, 295, 295, 296, 296, 297, 297, 298, 298, 303, 303, 304, 304, 305, 305, 306, 306, 311, 311, 312, 312, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 335, 335, 336, 336, 337, 337, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 345, 345, 346, 346, 359, 359, 360, 360, 361, 361, 362, 362, 363, 363, 364, 364, 365, 365, 366, 366, 383, 383, 384, 384, 385, 385, 386, 386, 387, 387, 388, 388, 389, 389, 390, 390, 391, 391, 392, 392, 393, 393, 394, 394, 395, 395, 396, 396, 397, 397, 398, 398, 447, 447, 448, 448, 449, 449, 450, 450, 451, 451, 452, 452, 453, 453, 454, 454, 455, 455, 456, 456, 457, 457, 458, 458, 459, 459, 460, 460, 461, 461, 462, 462),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 4, 4, 12, 12, 10, 10, 5, 5, 17, 17, 14, 14, 22, 22, 11, 11, 25, 25, 6, 6, 29, 29, 13, 13, 34, 34, 28, 28, 18, 18, 40, 40, 37, 37, 9, 9, 46, 46, 35, 35, 24, 24, 21, 21, 53, 53, 8, 8, 57, 57, 60, 60, 47, 47, 15, 15, 66, 66, 67, 67, 55, 55, 38, 38, 73, 73, 26, 26, 78, 78, 79, 79, 27, 27, 84, 84, 23, 23, 62, 62, 89, 89, 81, 81, 87, 87, 86, 86, 32, 32, 100, 100, 65, 65, 103, 103, 31, 31, 52, 52, 56, 56, 59, 59, 114, 114, 43, 43, 108, 108, 42, 42, 122, 122, 80, 80, 125, 125, 19, 19, 130, 130, 39, 39, 133, 133, 54, 54, 138, 138, 115, 115, 106, 106, 120, 120, 33, 33, 147, 147, 150, 150, 119, 119, 49, 49, 136, 136, 135, 135, 16, 16, 161, 161, 69, 69, 41, 41, 168, 168, 91, 91, 64, 64, 174, 174, 51, 51, 30, 30, 179, 179, 182, 182, 68, 68, 44, 44, 163, 163, 183, 183, 137, 137, 63, 63, 196, 196, 70, 70, 105, 105, 99, 99, 203, 203, 77, 77, 207, 207, 210, 210, 20, 20, 213, 213, 61, 61, 217, 217, 104, 104, 222, 222, 195, 195, 189, 189, 141, 141, 185, 185, 85, 85, 173, 173, 48, 48, 237, 237, 239, 239, 50, 50, 134, 134, 246, 246, 126, 126, 121, 121, 83, 83, 254, 254, 149, 149, 218, 218, 260, 260, 113, 113, 264, 264, 266, 266, 74, 74, 221, 221, 208, 208, 274, 274, 180, 180, 277, 277, 280, 280, 58, 58, 283, 283, 286, 286, 287, 287, 245, 245, 148, 148, 294, 294, 209, 209, 253, 253, 36, 36, 45, 45, 82, 82, 88, 88, 90, 90, 92, 92, 101, 101, 102, 102, 107, 107, 116, 116, 129, 129, 131, 131, 132, 132, 142, 142, 162, 162, 164, 164, 167, 167, 181, 181, 184, 184, 186, 186, 190, 190, 204, 204, 214, 214, 215, 215, 216, 216, 219, 219, 220, 220, 238, 238, 240, 240, 259, 259, 263, 263, 265, 265, 273, 273, 278, 278, 279, 279, 284, 284, 285, 285, 288, 288, 289, 289, 290, 290, 293, 293, 301, 301, 302, 302, 303, 303, 304, 304, 309, 309, 310, 310, 317, 317, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 329, 329, 330, 330, 331, 331, 332, 332, 335, 335, 336, 336, 345, 345, 346, 346, 355, 355, 356, 356, 361, 361, 362, 362, 367, 367, 368, 368, 371, 371, 372, 372, 373, 373, 374, 374, 375, 375, 376, 376, 387, 387, 388, 388, 389, 389, 390, 390, 407, 407, 408, 408, 409, 409, 410, 410, 435, 435, 436, 436, 437, 437, 438, 438, 439, 439, 440, 440, 441, 441, 442, 442, 447, 447, 448, 448, 449, 449, 450, 450, 451, 451, 452, 452, 453, 453, 454, 454, 463, 463, 464, 464, 465, 465, 466, 466, 467, 467, 468, 468, 469, 469, 470, 470),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 4, 4, 12, 12, 10, 10, 5, 5, 17, 17, 14, 14, 22, 22, 11, 11, 25, 25, 13, 13, 18, 18, 32, 32, 27, 27, 28, 28, 16, 16, 30, 30, 39, 39, 8, 8, 45, 45, 48, 48, 9, 9, 52, 52, 21, 21, 53, 53, 6, 6, 59, 59, 19, 19, 26, 26, 66, 66, 62, 62, 15, 15, 71, 71, 47, 47, 76, 76, 29, 29, 20, 20, 31, 31, 65, 65, 50, 50, 60, 60, 89, 89, 72, 72, 49, 49, 61, 61, 46, 46, 99, 99, 102, 102, 90, 90, 23, 23, 24, 24, 33, 33, 34, 34, 35, 35, 36, 36, 37, 37, 38, 38, 40, 40, 41, 41, 42, 42, 43, 43, 44, 44, 51, 51, 54, 54, 55, 55, 56, 56, 57, 57, 58, 58, 63, 63, 64, 64, 67, 67, 68, 68, 69, 69, 70, 70, 73, 73, 74, 74, 75, 75, 77, 77, 78, 78, 79, 79, 80, 80, 81, 81, 82, 82, 83, 83, 84, 84, 85, 85, 86, 86, 87, 87, 88, 88, 91, 91, 92, 92, 93, 93, 94, 94, 95, 95, 96, 96, 97, 97, 98, 98, 100, 100, 101, 101, 103, 103, 104, 104, 105, 105, 106, 106, 107, 107, 108, 108, 109, 109, 110, 110, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 117, 117, 118, 118, 119, 119, 120, 120, 121, 121, 122, 122, 123, 123, 124, 124, 125, 125, 126, 126, 127, 127, 128, 128, 129, 129, 130, 130, 131, 131, 132, 132, 133, 133, 134, 134, 135, 135, 136, 136, 137, 137, 138, 138, 139, 139, 140, 140, 141, 141, 142, 142, 143, 143, 144, 144, 145, 145, 146, 146, 147, 147, 148, 148, 149, 149, 150, 150, 151, 151, 152, 152, 153, 153, 154, 154, 155, 155, 156, 156, 157, 157, 158, 158, 159, 159, 160, 160, 161, 161, 162, 162, 163, 163, 164, 164, 165, 165, 166, 166, 167, 167, 168, 168, 169, 169, 170, 170, 171, 171, 172, 172, 173, 173, 174, 174, 175, 175, 176, 176, 177, 177, 178, 178, 179, 179, 180, 180, 181, 181, 182, 182, 183, 183, 184, 184, 185, 185, 186, 186, 187, 187, 188, 188, 189, 189, 190, 190, 191, 191, 192, 192, 193, 193, 194, 194, 195, 195, 196, 196, 197, 197, 198, 198, 199, 199, 200, 200, 201, 201, 202, 202, 203, 203, 204, 204, 205, 205, 206, 206, 207, 207, 208, 208, 209, 209, 210, 210, 211, 211, 212, 212, 213, 213, 214, 214, 247, 247, 248, 248, 249, 249, 250, 250, 267, 267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 272, 273, 273, 274, 274, 323, 323, 324, 324, 325, 325, 326, 326, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 412, 412, 413, 413, 414, 414, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446, 463, 463, 464, 464, 465, 465, 466, 466, 467, 467, 468, 468, 469, 469, 470, 470)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 6, 6, 5, 5, 5, 5, 6, 6, 5, 5, 6, 6, 6, 6, 7, 7, 6, 6, 5, 5, 7, 7, 6, 6, 7, 7, 7, 7, 6, 6, 6, 6, 8, 8, 6, 6, 7, 7, 7, 7, 7, 7, 4, 4, 5, 5, 6, 6, 6, 6, 6, 6, 8, 8, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 5, 5, 6, 6, 8, 8, 7, 7, 7, 7, 8, 8, 7, 7, 3, 3, 4, 4, 8, 8, 8, 8, 8, 8, 5, 5, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 8, 8, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 5, 5, 8, 8, 5, 5, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 6, 6, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 6, 6, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 5, 5, 5, 5, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 5, 5, 6, 6, 7, 7, 4, 4, 5, 5, 7, 7, 7, 7, 6, 6, 7, 7, 3, 3, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 6, 6, 8, 8, 8, 8, 5, 5, 6, 6, 8, 8, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 5, 5, 6, 6, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 5, 5, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 4, 4, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 5, 5, 6, 6, 6, 6, 3, 3, 4, 4, 5, 5, 4, 4, 5, 5, 6, 6, 6, 6, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 6, 6, 5, 5, 6, 6, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 4, 4, 5, 5, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((61, 62, 81, 82, 89, 90, 91, 92, 101, 102, 107, 108, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126, 127, 128, 131, 132, 135, 136, 139, 140, 141, 142, 147, 148, 149, 150, 151, 152, 157, 158, 159, 160, 167, 168, 173, 174, 177, 178, 179, 180, 181, 182, 183, 184, 189, 190, 191, 192, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 213, 214, 215, 216, 221, 222, 229, 230, 231, 232, 237, 238, 239, 240, 249, 250, 253, 254, 255, 256, 259, 260, 261, 262, 263, 264, 271, 272, 275, 276, 277, 278, 279, 280, 281, 282, 287, 288, 289, 290, 299, 300, 301, 302, 307, 308, 309, 310, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510),
                (71, 72, 75, 76, 93, 94, 95, 96, 97, 98, 109, 110, 111, 112, 117, 118, 123, 124, 127, 128, 139, 140, 143, 144, 145, 146, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 165, 166, 169, 170, 171, 172, 175, 176, 177, 178, 187, 188, 191, 192, 193, 194, 197, 198, 199, 200, 201, 202, 205, 206, 211, 212, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 241, 242, 243, 244, 247, 248, 249, 250, 251, 252, 255, 256, 257, 258, 261, 262, 267, 268, 269, 270, 271, 272, 275, 276, 281, 282, 291, 292, 295, 296, 297, 298, 299, 300, 305, 306, 307, 308, 311, 312, 313, 314, 315, 316, 323, 324, 325, 326, 327, 328, 333, 334, 337, 338, 339, 340, 341, 342, 343, 344, 347, 348, 349, 350, 351, 352, 353, 354, 357, 358, 359, 360, 363, 364, 365, 366, 369, 370, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 443, 444, 445, 446, 455, 456, 457, 458, 459, 460, 461, 462, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510),
                (215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
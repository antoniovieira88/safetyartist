library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 1, 2, 0, 0, 1, 1, 1, 2, 1, 2, 1, 0, 0, 0, 2, 2, 0, 2, 2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 1, 2, 0, 1, -2, -2, 0, 2, 1, 0, -2, 2, -2, 1, 0, 1, 0, -2, 0, -2, 1, 2, -2, 2, 2, 1, 1, 2, -2, 0, -2, 1, 1, 1, -2, 0, 2, 1, 0, 0, 1, 1, 1, 1, 1, -2, 0, 1, 2, 1, 1, 2, 0, 0, -2, 1, 1, 0, -2, 2, 1, 1, -2, -2, 0, 2, -2, 1, 1, -2, 0, 0, -2, -2, 1, -2, 2, -2, -2, -2, 0, -2, 1, 1, -2, 1, 1, 1, -2, 0, -2, 2, -2, -2, -2, 0, 1, -2, -2, -2, 2, -2, 2, 0, -2, -2, -2, -2, 1, 1, -2, -2, -2, -2, 1, 0, -2, -2, 2, -2, 1, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 0, 2, -2, -2, -2, -2, -2, 0, 0, 2, 0, 0, 2, 0, -2, 0, 0, -2, 0, -2, -2, -2, -2, -2, -2, 1, 2, 0, 0, -2, 1, 0, 1, 1, 0, -2, -2, 1, -2, 0, -2, -2, -2, -2, 0, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 1, 1, 2, 1, -2, 2, -2, -2, -2, -2, 1, 1, -2, 2, -2, -2, -2, 0, -2, -2, -2, 1, 2, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, 0, -2, -2, 1, -2, 1, -2, -2, -2, -2, -2, -2, 1, 2, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, 1, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, 1, 0, -2, -2, 2, -2, -2, -2, 2, -2, -2, -2, -2, 0, -2, -2, -2, 2, 0, -2, 1, -2, -2, -2, -2, 1, -2, -2, 1, 1, -2, 2, -2, -2, 1, -2, -2, -2, -2, -2, -2, 0, 2, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 1, 2, 1, 0, 0, 1, 1, 2, 2, 0, 0, 1, 1, 1, 2, 1, 0, 1, 2, 2, 0, 0, 0, 2, 0, 1, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, -2, 0, 1, 0, 2, 0, 0, -2, 1, 1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, -2, 1, 0, 2, -2, 2, 1, 1, 1, 0, 1, 2, 1, 1, -2, 0, 2, 0, 1, 1, 1, 1, -2, -2, 0, 1, -2, 0, -2, -2, 0, 0, 1, 2, 0, -2, 1, 1, 0, -2, 1, 0, 0, 0, 2, 0, -2, -2, -2, -2, -2, 2, -2, 1, -2, -2, 1, 2, -2, -2, 1, 2, -2, 0, 1, 0, -2, 2, 0, -2, 0, 2, -2, 1, -2, -2, 1, 0, 1, 2, 0, 2, -2, -2, 0, 1, 0, 2, -2, -2, 2, 2, 1, 1, -2, 0, -2, -2, -2, 0, 2, 2, -2, -2, 0, 1, 0, 0, -2, -2, 0, 1, 0, 1, 1, -2, -2, 1, 2, 1, 0, 2, 1, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, 1, -2, -2, 1, -2, -2, 1, 1, -2, -2, -2, -2, -2, -2, -2, 1, 0, 0, -2, -2, 0, 1, 2, -2, 1, 1, -2, 2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, 1, 2, -2, -2, 0, 0, -2, -2, -2, -2, 1, -2, -2, 1, 1, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 0, -2, 1, -2, -2, -2, 1, 1, 1, 2, -2, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, 2, -2, 1, -2, -2, 1, -2, 1, 1, -2, -2, -2, -2, 2, 0, -2, -2, -2, -2, 2, 0, -2, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, 2, 0, -2, 0, 1, -2, -2, -2, -2, -2, -2, -2, 2, 0, -2, -2, -2, -2, 0, -2, -2, -2, 0, 1, 1, -2, -2, 0, -2, -2, 2, -2, -2, -2, -2, -2, -2, 0, 1, -2, 1, 2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, -2, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((1145163, 55893, 1806227, 277007, 820053, 22073, 40953, 85844, 2283949, 76119, 4285, 76573, 29734, 96666, 101403, 65094, 75228, 3502, 89293, 6029, 117653, 329060, 486055, 418114, 619596, 1303922, 1565176, 1360628, 5238, 63401, 4285, 884077, 1027253, 73895, 2929, 1510150, 1393618, 97697, 109638, 94146, 3502, 106724, 4285, 76948, 1713617, 1587665, 1675876, 3502, 2929, 1765031, 3502, 4285, -8192, 1124693, 984207, 86240, 83906, 172705, 245934, 164602, 214447, 656075, 694414, 582148, 3502, 57449, 4285, 3502, 2929, 46962, 4285, 20361, 7032, -8192, -8192, 534851, 2929, 97877, 1351029, -8192, 5238, -8192, 114720, 976992, 70665, 1058458, -8192, 2051331, -8192, 45663, 3502, -8192, 4285, 3502, 85432, 78140, 4285, -8192, 1394286, -8192, 92387, 13251, 18054, -8192, 86893, 2929, 107549, 2247623, 2007933, 101916, 104261, 111648, 114239, 105173, -8192, 1293759, 80186, 5238, 99294, 86791, 2929, 2071333, 1843500, -8192, 95659, 31408, 372572, -8192, 4285, 34959, 37824, -8192, -8192, 499512, 4285, -8192, 61512, 111387, -8192, 1679603, 1664326, -8192, -8192, 99898, -8192, 5238, -8192, -8192, -8192, 903631, -8192, 64764, 72311, -8192, 67479, 59532, 64897, -8192, 764030, -8192, 5238, -8192, -8192, -8192, 811413, 82519, -8192, -8192, -8192, 5238, -8192, 4285, 328842, -8192, -8192, -8192, -8192, 88899, 96688, -8192, -8192, -8192, -8192, 50180, 493637, -8192, -8192, 4285, -8192, 27833, -8192, -8192, -8192, 59295, 1006085, -8192, -8192, -8192, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, -8192, 93852, -8192, -8192, -8192, -8192, 142783, 4285, -8192, -8192, -8192, -8192, -8192, 2344752, 2743214, 2929, 2868247, 2617507, 3502, 2335336, -8192, 2302480, 2404686, -8192, 1034935, -8192, -8192, -8192, -8192, -8192, -8192, 69565, 2929, 1368785, 1225857, -8192, 75132, 740952, 55824, 50822, 773430, -8192, -8192, 82551, -8192, 1573908, -8192, -8192, -8192, -8192, 2130333, -8192, -8192, -8192, -8192, 44596, -8192, -8192, -8192, -8192, -8192, 68555, 70172, 4285, 79091, -8192, 5238, -8192, -8192, -8192, -8192, 96343, 100116, -8192, 5238, -8192, -8192, -8192, 2701964, -8192, -8192, -8192, 102246, 3502, 104050, -8192, 99811, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 5238, -8192, -8192, 746171, -8192, -8192, 37569, -8192, 35855, -8192, -8192, -8192, -8192, -8192, -8192, 35083, 4285, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 5238, -8192, 59372, -8192, -8192, -8192, -8192, -8192, -8192, 945420, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 1184907, 70457, 1277553, -8192, -8192, 2929, -8192, -8192, -8192, 2929, -8192, -8192, -8192, -8192, 1139332, -8192, -8192, -8192, 2929, 1923317, -8192, 89133, -8192, -8192, -8192, -8192, 100307, -8192, -8192, 100955, 105987, -8192, 2929, -8192, -8192, 103453, -8192, -8192, -8192, -8192, -8192, -8192, 2623701, 2929, -8192, 107214, -8192, -8192, -8192, 68500, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192),
                (1396964, 52341, 2049265, 360371, 867137, 24262, 498698, 89907, 2375670, 81132, 4285, 99491, 106549, 61793, 70824, 2929, 85422, 121294, 255447, 8402, 18223, 4285, 5238, 1308907, 991861, 41507, 49603, 38102, 4285, 101917, 2705376, 96719, 3502, 2929, 2098257, 1432907, 1750936, 5238, 1768288, 77524, 2929, 1844013, 3502, 3502, 1926221, 1849363, 1675978, 1697507, 1885490, 614799, 739112, 499989, 4285, 731681, 633773, 93865, -8192, 1716529, 115136, 1074079, 2929, 21345, 79886, -8192, 7062, 27565, 34299, 32374, 5238, 77153, 1071550, 4285, 96076, 1034347, 1353086, 86855, 1138092, 65931, 977378, 981968, 1166462, -8192, 69034, 726826, 3502, -8192, 5238, 42934, 45838, 44863, 409746, 94250, 2929, 54704, 60009, -8192, 156412, 4285, 184353, 75235, 79365, 92622, 97721, -8192, -8192, 1231576, 103038, -8192, 61804, -8192, -8192, 1490305, 1558582, 92906, 2929, 2230636, -8192, 57610, 65333, 1564138, -8192, 86909, 1662086, 571872, 608840, 3502, 735605, -8192, -8192, -8192, -8192, -8192, 4285, -8192, 62455, -8192, -8192, 71172, 3502, -8192, -8192, 33462, 2929, -8192, 370654, 65396, 1024691, -8192, 4285, 925531, -8192, 492178, 4285, -8192, 55846, -8192, -8192, 105762, 2887680, 102253, 2929, 2546238, 3502, -8192, -8192, 1553068, 97241, 533653, 5238, -8192, -8192, 3502, 3502, 101008, 105352, -8192, 2043439, -8192, -8192, -8192, 1564634, 2929, 2929, -8192, -8192, 1396425, 92539, 1181538, 1374904, -8192, -8192, 185582, 31924, 162618, 26332, 25317, -8192, -8192, 13059, 4285, 15486, 284186, 3502, 37105, 40116, -8192, 43595, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 2929, -8192, 50794, -8192, -8192, 50793, -8192, -8192, 82663, 85259, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 106144, 2230089, 2371572, -8192, -8192, 692239, 76002, 4285, -8192, 66524, 69889, -8192, 5238, -8192, -8192, -8192, -8192, -8192, -8192, 1493308, -8192, -8192, -8192, 102747, -8192, 101529, 5238, -8192, -8192, 454241, 482798, -8192, -8192, -8192, -8192, 107533, -8192, -8192, 98994, 86245, -8192, -8192, -8192, -8192, -8192, 80565, -8192, -8192, -8192, -8192, -8192, 2479187, -8192, 111746, -8192, -8192, -8192, 45994, 47781, 43732, 2929, -8192, 538046, 4285, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 1766896, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 4285, -8192, -8192, 4285, -8192, 110969, -8192, -8192, 114002, -8192, 112843, 111036, -8192, -8192, -8192, -8192, 2929, 393280, -8192, -8192, -8192, -8192, 2929, 2591141, -8192, 104350, -8192, 29336, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 1535835, -8192, -8192, -8192, -8192, -8192, 112902, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 690380, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 100669, -8192, -8192, -8192, -8192, -8192, 66903, -8192, -8192, -8192, 109473, -8192, -8192, 2929, 2788154, -8192, 2748997, 111775, -8192, -8192, -8192, -8192, -8192, -8192, -8192, 2929, 1555822, -8192, -8192, -8192, -8192, 494478, -8192, -8192, -8192, 1801411, 101593, 105749, -8192, -8192, 204101, -8192, -8192, 3502, -8192, -8192, -8192, -8192, -8192, -8192, 650206, 63346, -8192, 67665, 4285, -8192, -8192, -8192, -8192, 46347, -8192, -8192, -8192, -8192, 66293, -8192, -8192, -8192, -8192, 93342, -8192, -8192, -8192, 47878, -8192, -8192, -8192, 650383, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192),
                (2082780, 53336, 2866606, 542776, 1187550, -8192, -8192, -8192, -8192, 99874, 2874724, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192, -8192)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((1228, 586, 1334, 1054, 139, 444, 1256, 1107, 1357, 1331, 445, 953, 96, 139, 915, 37, 412, 1045, 114, 223, 1251, 1348, 1002, 195, 1262, 1242, 530, 237, 1142, 689, 1279, 1220, 310, 1359, 1092, 546, 1232, 1276, 1364, 1354, 832, 228, 1254, 43, 1122, 382, 21, 145, 832, 124, 1203, 327, 0, 11, 785, 434, 1143, 369, 12, 18, 1131, 185, 9, 48, 788, 202, 1148, 1001, 1336, 554, 1245, 708, 21, 0, 1365, 1170, 178, 803, 1332, 0, 506, 0, 975, 65, 740, 1268, 0, 1000, 1365, 81, 569, 0, 1205, 1035, 1356, 416, 1245, 0, 467, 0, 986, 931, 1328, 1365, 91, 390, 19, 111, 715, 303, 1024, 755, 1283, 989, 0, 1138, 161, 998, 171, 1363, 1143, 431, 1345, 0, 1024, 1183, 1361, 1365, 592, 216, 1241, 1260, 273, 14, 364, 0, 993, 874, 1365, 1195, 303, 1092, 0, 31, 819, 579, 0, 303, 910, 1097, 1365, 683, 1293, 1365, 137, 819, 1318, 1365, 341, 1365, 887, 341, 1252, 819, 62, 975, 1365, 1365, 341, 281, 0, 105, 853, 0, 1365, 1365, 546, 735, 1260, 1365, 455, 1260, 768, 986, 1338, 1365, 512, 934, 1365, 546, 1365, 910, 0, 780, 1297, 1365, 341, 0, 910, 455, 1365, 585, 0, 0, 1024, 1195, 683, 1006, 1365, 1268, 273, 1365, 1145, 390, 1365, 0, 910, 0, 546, 1365, 1339, 1053, 1363, 105, 1287, 1062, 1365, 228, 1300, 1365, 910, 455, 1365, 0, 683, 0, 410, 1363, 1241, 910, 1339, 0, 1241, 1234, 1361, 780, 1342, 1365, 195, 986, 1365, 1155, 546, 819, 1365, 1365, 975, 455, 1365, 455, 0, 910, 1365, 1365, 455, 0, 390, 1, 54, 420, 20, 0, 1092, 819, 1365, 910, 1365, 1161, 1356, 1365, 853, 0, 1365, 0, 341, 683, 0, 0, 99, 341, 22, 0, 1138, 390, 0, 975, 1365, 910, 1365, 0, 273, 0, 683, 1365, 910, 0, 455, 910, 1365, 114, 0, 0, 546, 0, 1092, 1287, 1365, 1349, 0, 1365, 910, 0, 455, 0, 132, 683, 0, 0, 1365, 910, 1365, 1365, 910, 1248, 1365, 546, 1365, 1365, 1024, 1365, 910, 910, 1365, 455, 0, 0, 111, 0, 683, 0, 455, 1365, 1092, 0, 273, 1170, 1365, 1365, 910, 273, 0, 1092, 1365, 1092, 1365, 1092, 1365, 273, 0, 1365, 910, 455, 0, 910, 455, 910, 1365, 1365, 1323, 956, 1347, 0, 1365, 1214, 1365, 819, 1365, 195, 0, 0, 455, 0, 171, 455, 0, 1365, 1331, 1183, 1365, 585, 1365, 910, 341, 1365, 1260, 910, 1365, 1349, 1365, 1365, 1145, 0, 1365, 98, 0, 0, 455, 105, 0, 1365, 1359, 1203, 1365, 228, 1365, 0, 455, 10, 0, 0, 455, 0, 0, 0, 0, 1365, 1365, 0, 0, 0, 0, 0, 0, 1365, 1365, 0, 0, 0, 0, 0, 0, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 819, 819, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 819, 819, 1365, 1365, 0, 0, 1365, 1365, 546, 546, 1365, 1365, 1365, 1365, 1365, 1365, 341, 341, 455, 455, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 546, 546, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 546, 546, 1365, 1365, 1365, 1365, 0, 0, 819, 819, 1365, 1365, 1365, 1365, 0, 0, 683, 683, 0, 0, 0, 0, 0, 0, 910, 910, 1365, 1365, 0, 0, 1365, 1365, 910, 910, 0, 0, 455, 455, 0, 0, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 910, 910, 0, 0, 455, 455, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 546, 546, 1365, 1365, 1365, 1365, 1024, 1024, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 0, 0, 0, 0, 0, 0, 455, 455, 1365, 1365, 1092, 1092, 0, 0, 273, 273, 1365, 1365, 273, 273, 0, 0, 1092, 1092, 1365, 1365, 273, 273, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 455, 455, 0, 0, 455, 455, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 455, 455, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 819, 819, 819, 819, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 546, 546, 546, 546, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1092, 1092, 1092, 1092, 0, 0, 0, 0, 273, 273, 273, 273, 273, 273, 273, 273, 0, 0, 0, 0, 1092, 1092, 1092, 1092, 1365, 1365, 1365, 1365, 273, 273, 273, 273, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 455, 455, 455, 455, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
                (1093, 409, 1321, 932, 138, 320, 1286, 1045, 1355, 1331, 405, 153, 1044, 31, 368, 1219, 176, 734, 85, 220, 1254, 476, 68, 189, 1145, 966, 1347, 1310, 237, 1234, 1362, 1349, 610, 90, 1328, 1291, 730, 396, 1339, 1364, 1060, 435, 1267, 384, 46, 187, 898, 158, 1285, 174, 9, 38, 656, 361, 1336, 443, 1365, 72, 910, 109, 711, 566, 61, 0, 1105, 26, 330, 1161, 89, 666, 1317, 26, 278, 732, 95, 171, 1218, 890, 1303, 1134, 410, 0, 1229, 53, 657, 1365, 341, 76, 627, 1274, 186, 75, 559, 406, 1205, 1365, 1011, 171, 1218, 273, 1024, 253, 1044, 1195, 188, 35, 683, 1365, 585, 0, 1365, 1155, 273, 1364, 1102, 216, 1365, 683, 1332, 1045, 1365, 341, 1280, 1359, 1173, 359, 1306, 1365, 569, 1365, 273, 0, 975, 1365, 341, 853, 0, 8, 232, 101, 662, 1343, 887, 0, 1183, 1096, 1356, 1365, 768, 410, 1365, 3, 230, 0, 735, 910, 0, 1318, 1365, 1362, 905, 103, 1302, 1365, 372, 840, 228, 1214, 482, 0, 910, 12, 203, 19, 683, 1365, 241, 137, 853, 546, 1312, 883, 1337, 0, 1155, 1, 110, 432, 19, 64, 1365, 193, 6, 21, 975, 455, 1365, 0, 280, 1170, 85, 1280, 683, 35, 390, 1365, 161, 512, 1365, 0, 1092, 819, 1365, 759, 1365, 1006, 1365, 228, 1365, 0, 683, 455, 1365, 65, 546, 1365, 0, 910, 94, 0, 910, 0, 217, 637, 85, 0, 1365, 2, 58, 306, 0, 16, 1101, 1365, 853, 228, 1229, 98, 910, 137, 683, 607, 0, 228, 1365, 1162, 1365, 1327, 621, 195, 1365, 341, 18, 0, 1365, 910, 0, 26, 546, 0, 512, 993, 1365, 1365, 546, 420, 0, 1128, 1365, 1365, 759, 0, 546, 1158, 1365, 745, 1365, 1092, 455, 1281, 1365, 1342, 683, 0, 1024, 241, 0, 98, 910, 390, 0, 1365, 910, 455, 0, 683, 1365, 146, 0, 99, 683, 910, 273, 0, 171, 512, 0, 1365, 1092, 455, 1365, 1170, 1365, 910, 1365, 1365, 683, 0, 218, 420, 0, 273, 910, 1365, 1229, 585, 1365, 0, 1024, 1365, 1252, 910, 1365, 585, 1365, 1062, 1365, 1365, 455, 455, 0, 910, 1365, 819, 1365, 341, 910, 910, 1365, 7, 210, 248, 0, 0, 910, 0, 341, 61, 455, 0, 341, 1365, 910, 910, 1365, 273, 0, 28, 341, 910, 1365, 1365, 1024, 1092, 1365, 1365, 1092, 455, 910, 455, 0, 455, 910, 228, 0, 0, 455, 1365, 1138, 1271, 1365, 1365, 455, 1351, 1365, 1365, 1146, 643, 1365, 228, 869, 1092, 683, 0, 455, 119, 0, 1365, 1329, 1179, 1365, 546, 1365, 0, 105, 455, 0, 0, 37, 11, 152, 585, 0, 38, 0, 0, 241, 0, 683, 1241, 1365, 91, 0, 0, 21, 683, 11, 171, 0, 0, 910, 0, 85, 455, 0, 0, 76, 62, 0, 0, 455, 1365, 1330, 910, 1365, 1365, 1343, 910, 1365, 0, 6, 455, 0, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 1365, 1365, 546, 546, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1092, 1092, 1365, 1365, 1365, 1365, 0, 0, 455, 455, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 0, 0, 1365, 1365, 546, 546, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 546, 546, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 683, 683, 1365, 1365, 0, 0, 910, 910, 273, 273, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 0, 0, 341, 341, 455, 455, 0, 0, 341, 341, 1365, 1365, 910, 910, 341, 341, 1365, 1365, 1024, 1024, 1092, 1092, 1365, 1365, 1365, 1365, 1092, 1092, 0, 0, 1365, 1365, 1365, 1365, 455, 455, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 546, 546, 1365, 1365, 0, 0, 455, 455, 0, 0, 0, 0, 0, 0, 0, 0, 683, 683, 0, 0, 0, 0, 0, 0, 1365, 1365, 910, 910, 1365, 1365, 1365, 1365, 910, 910, 1365, 1365, 0, 0, 455, 455, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 546, 546, 546, 546, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 1092, 1092, 1092, 1092, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 546, 546, 546, 546, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 683, 683, 683, 683, 1365, 1365, 1365, 1365, 910, 910, 910, 910, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 546, 546, 546, 546, 546, 546, 546, 546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365),
                (682, 208, 1329, 623, 87, 176, 1335, 21, 304, 1132, 1365, 1355, 522, 1339, 1365, 176, 176, 1335, 1335, 21, 21, 304, 304, 1355, 1355, 522, 522, 1339, 1339, 1365, 1365, 176, 176, 176, 176, 1335, 1335, 1335, 1335, 21, 21, 21, 21, 304, 304, 304, 304, 1355, 1355, 1355, 1355, 522, 522, 522, 522, 1339, 1339, 1339, 1339, 1365, 1365, 1365, 1365, 176, 176, 176, 176, 176, 176, 176, 176, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 21, 21, 21, 21, 21, 21, 21, 21, 304, 304, 304, 304, 304, 304, 304, 304, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 522, 522, 522, 522, 522, 522, 522, 522, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 1335, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 304, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 1355, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 522, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1339, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365, 1365)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 7, 5, 15, 11, 21, 9, 37, 33, 13, 19, 57, 45, 25, 61, 17, 29, 51, 71, 101, 125, 23, 89, 67, 77, 27, 79, 137, 31, 149, 193, 83, 237, 35, 43, 93, 39, 219, 119, 41, 105, 87, 367, 249, 47, 287, 97, 49, 217, 207, 53, 431, 391, 55, 145, 159, 59, 323, 353, 187, 63, 267, 133, 65, 163, 155, 69, 243, 75, 183, 73, 359, 433, 435, 275, 235, 117, 277, 437, 81, 439, 141, 299, 85, 329, 441, 111, 443, 169, 91, 445, 261, 95, 351, 115, 165, 447, 99, 449, 131, 103, 211, 451, 321, 107, 387, 143, 109, 259, 205, 113, 255, 181, 453, 375, 293, 177, 349, 395, 121, 123, 297, 455, 199, 127, 315, 457, 129, 201, 339, -1, -1, 345, 135, 459, 175, 139, 461, 295, 233, -1, -1, 417, 463, 147, 465, -1, -1, 151, 467, 153, 229, 469, 343, 157, 303, 471, 197, 473, 161, -1, -1, 475, 305, 167, 477, -1, -1, 171, 479, 265, 173, -1, -1, 481, 483, 179, 331, -1, -1, -1, -1, 185, 365, -1, -1, 189, 485, 191, 487, -1, -1, 195, 355, 489, 491, -1, -1, 493, 495, 203, 497, -1, -1, -1, -1, 209, 499, -1, -1, 501, 213, 215, 503, -1, -1, 505, 507, 407, 221, 223, 333, 283, 225, 227, 509, 371, 307, 511, 231, -1, -1, -1, -1, -1, -1, 377, 239, 241, 363, 513, 341, 245, 337, 247, 361, -1, -1, 251, 515, 253, 517, -1, -1, 519, 257, -1, -1, -1, -1, 263, 521, -1, -1, -1, -1, 427, 269, 271, 309, 523, 273, 525, 527, -1, -1, 279, 403, 529, 281, -1, -1, 531, 285, 533, 535, 537, 289, 291, 413, 539, 369, -1, -1, -1, -1, 541, 543, 545, 301, -1, -1, 547, 549, 551, 553, -1, -1, 311, 555, 557, 313, -1, -1, 317, 559, 319, 561, 563, 565, 567, 569, 571, 325, 327, 573, 575, 577, -1, -1, -1, -1, 335, 579, 581, 583, 585, 587, 589, 591, 593, 595, -1, -1, 597, 347, 599, 373, 601, 603, 605, 607, 609, 611, 357, 613, -1, -1, 615, 617, -1, -1, 619, 621, -1, -1, 623, 625, -1, -1, -1, -1, -1, -1, -1, -1, 627, 379, 381, 383, 629, 631, 385, 633, -1, -1, 389, 635, 637, 639, 641, 393, 643, 645, 647, 397, 399, 649, 401, 651, -1, -1, 653, 405, -1, -1, 409, 419, 655, 411, 657, 659, 415, 661, -1, -1, -1, -1, 663, 421, 423, 665, 425, 667, -1, -1, 429, 669, 671, 673, 675, 677, 679, 681, 683, 685, 687, 689, -1, -1, -1, -1, 691, 693, 695, 697, 699, 701, -1, -1, 703, 705, -1, -1, 707, 709, 711, 713, 715, 717, 719, 721, -1, -1, -1, -1, 723, 725, -1, -1, -1, -1, -1, -1, 727, 729, -1, -1, 731, 733, -1, -1, -1, -1, 735, 737, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 739, 741, -1, -1, -1, -1, -1, -1, 743, 745, -1, -1, 747, 749, 751, 753, -1, -1, -1, -1, -1, -1, 755, 757, -1, -1, -1, -1, -1, -1, 759, 761, -1, -1, -1, -1, 763, 765, -1, -1, 767, 769, 771, 773, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 775, 777, -1, -1, 779, 781, 783, 785, -1, -1, -1, -1, -1, -1, -1, -1, 787, 789, 791, 793, -1, -1, -1, -1, 795, 797, 799, 801, 803, 805, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 807, 809, -1, -1, -1, -1, -1, -1, 811, 813, 815, 817, 819, 821, 823, 825, -1, -1, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, 847, 849, 851, 853, -1, -1, -1, -1, -1, -1, 855, 857, -1, -1, -1, -1, 859, 861, -1, -1, -1, -1, 863, 865, 867, 869, -1, -1, -1, -1, 871, 873, 875, 877, 879, 881, -1, -1, 883, 885, 887, 889, -1, -1, 891, 893, 895, 897, 899, 901, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, 951, 953, 955, 957, -1, -1, -1, -1, 959, 961, 963, 965, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, -1, -1, -1, -1, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, -1, -1, -1, -1, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 13, 17, 25, 9, 29, 39, 11, 43, 35, 49, 15, 77, 21, 19, 65, 61, 95, 23, 71, 59, 69, 27, 123, 141, 87, 31, 157, 113, 33, 231, 321, 179, 37, 57, 351, 417, 41, 47, 119, 45, 171, 91, 55, 223, 357, 51, 237, 151, 53, 83, 383, 165, 473, 267, 111, 137, 99, 63, 197, 475, 107, 191, 67, 201, 203, 85, 277, 185, 73, 75, 105, 227, 211, 79, 145, 117, 81, 477, 371, 377, 93, 479, 177, 261, 89, 381, 219, 307, 101, 103, 301, 481, 97, 281, 181, 155, 127, 135, 129, -1, -1, 313, 163, 483, 109, -1, -1, 213, 229, 461, 115, 269, 485, 133, 385, 121, 487, 251, 271, 289, 125, 131, 215, -1, -1, -1, -1, 489, 305, 491, 315, -1, -1, 375, 139, -1, -1, 333, 143, 493, 221, 147, 399, 495, 149, 249, 497, 423, 153, 499, 167, -1, -1, 159, 403, 339, 161, 327, 283, -1, -1, 207, 275, 373, 169, -1, -1, 427, 173, 393, 175, 501, 247, -1, -1, 503, 255, 183, 439, -1, -1, 365, 187, 189, 359, -1, -1, 193, 433, 369, 195, 265, 505, 507, 199, 379, 299, 345, 209, 295, 205, 509, 303, -1, -1, 511, 513, -1, -1, -1, -1, 217, 515, 389, 517, 519, 391, 521, 523, 361, 225, 525, 527, -1, -1, -1, -1, 529, 233, 235, 367, 531, 533, 443, 239, 241, 535, 457, 243, 537, 245, -1, -1, -1, -1, -1, -1, 253, 539, -1, -1, 257, 541, 397, 259, -1, -1, 263, 451, 543, 545, -1, -1, 349, 547, 549, 311, 273, 551, -1, -1, -1, -1, 279, 553, -1, -1, 555, 557, 285, 559, 287, 561, -1, -1, 291, 465, 317, 293, 563, 353, 297, 565, -1, -1, -1, -1, -1, -1, -1, -1, 567, 569, 309, 571, -1, -1, 573, 575, -1, -1, -1, -1, 577, 319, -1, -1, 323, 579, 325, 581, 583, 387, 585, 329, 331, 587, -1, -1, 589, 335, 337, 591, -1, -1, 593, 341, 343, 595, 355, 597, 347, 599, -1, -1, -1, -1, 601, 603, -1, -1, -1, -1, 605, 607, -1, -1, 363, 609, -1, -1, 611, 613, 415, 615, 617, 619, 621, 623, -1, -1, -1, -1, 455, 625, -1, -1, 627, 629, 631, 633, 635, 637, -1, -1, -1, -1, -1, -1, 395, 639, -1, -1, -1, -1, 401, 641, 643, 645, 405, 647, 649, 407, 409, 651, 413, 411, -1, -1, -1, -1, -1, -1, 653, 419, 421, 655, 657, 659, 661, 425, 663, 665, 667, 429, 441, 431, -1, -1, 435, 669, 671, 437, -1, -1, -1, -1, -1, -1, 469, 445, 673, 447, 449, 675, -1, -1, 677, 453, -1, -1, -1, -1, 459, 679, -1, -1, 681, 463, 683, 685, 687, 467, 689, 691, 693, 471, 695, 697, 699, 701, 703, 705, 707, 709, -1, -1, 711, 713, -1, -1, 715, 717, 719, 721, 723, 725, -1, -1, 727, 729, 731, 733, -1, -1, 735, 737, -1, -1, 739, 741, -1, -1, 743, 745, -1, -1, -1, -1, -1, -1, 747, 749, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 751, 753, -1, -1, -1, -1, 755, 757, -1, -1, -1, -1, 759, 761, -1, -1, -1, -1, -1, -1, 763, 765, -1, -1, -1, -1, -1, -1, -1, -1, 767, 769, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 771, 773, 775, 777, -1, -1, 779, 781, -1, -1, 783, 785, -1, -1, 787, 789, 791, 793, -1, -1, -1, -1, 795, 797, 799, 801, 803, 805, 807, 809, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 811, 813, 815, 817, -1, -1, -1, -1, -1, -1, 819, 821, -1, -1, -1, -1, 823, 825, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, 847, 849, 851, 853, -1, -1, -1, -1, 855, 857, 859, 861, -1, -1, 863, 865, -1, -1, -1, -1, -1, -1, 867, 869, 871, 873, 875, 877, 879, 881, -1, -1, -1, -1, 883, 885, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 887, 889, 891, 893, 895, 897, 899, 901, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 951, 953, 955, 957, 959, 961, 963, 965, -1, -1, -1, -1, 967, 969, 971, 973, 975, 977, 979, 981, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, 15, 17, 19, 21, 11, 13, 23, 25, 27, 29, 31, 33, 35, 37, 39, 41, 43, 45, 47, 49, 51, 53, 55, 57, 59, 61, 63, 65, 67, 69, 71, 73, 75, 77, 79, 81, 83, 85, 87, 89, 91, 93, 95, 97, 99, 101, 103, 105, 107, 109, 111, 113, 115, 117, 119, 121, 123, 125, 127, 129, 131, 133, 135, 137, 139, 141, 143, 145, 147, 149, 151, 153, 155, 157, 159, 161, 163, 165, 167, 169, 171, 173, 175, 177, 179, 181, 183, 185, 187, 189, 191, 193, 195, 197, 199, 201, 203, 205, 207, 209, 211, 213, 215, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 237, 239, 241, 243, 245, 247, 249, 251, 253, 255, 257, 259, 261, 263, 265, 267, 269, 271, 273, 275, 277, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 341, 343, 345, 347, 349, 351, 353, 355, 357, 359, 361, 363, 365, 367, 369, 371, 373, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 415, 417, 419, 421, 423, 425, 427, 429, 431, 433, 435, 437, 439, 441, 443, 445, 447, 449, 451, 453, 455, 457, 459, 461, 463, 465, 467, 469, 471, 473, 475, 477, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, 511, 513, 515, 517, 519, 521, 523, 525, 527, 529, 531, 533, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 555, 557, 559, 561, 563, 565, 567, 569, 571, 573, 575, 577, 579, 581, 583, 585, 587, 589, 591, 593, 595, 597, 599, 601, 603, 605, 607, 609, 611, 613, 615, 617, 619, 621, 623, 625, 627, 629, 631, 633, 635, 637, 639, 641, 643, 645, 647, 649, 651, 653, 655, 657, 659, 661, 663, 665, 667, 669, 671, 673, 675, 677, 679, 681, 683, 685, 687, 689, 691, 693, 695, 697, 699, 701, 703, 705, 707, 709, 711, 713, 715, 717, 719, 721, 723, 725, 727, 729, 731, 733, 735, 737, 739, 741, 743, 745, 747, 749, 751, 753, 755, 757, 759, 761, 763, 765, 767, 769, 771, 773, 775, 777, 779, 781, 783, 785, 787, 789, 791, 793, 795, 797, 799, 801, 803, 805, 807, 809, 811, 813, 815, 817, 819, 821, 823, 825, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, 847, 849, 851, 853, 855, 857, 859, 861, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, 887, 889, 891, 893, 895, 897, 899, 901, 903, 905, 907, 909, 911, 913, 915, 917, 919, 921, 923, 925, 927, 929, 931, 933, 935, 937, 939, 941, 943, 945, 947, 949, 951, 953, 955, 957, 959, 961, 963, 965, 967, 969, 971, 973, 975, 977, 979, 981, 983, 985, 987, 989, 991, 993, 995, 997, 999, 1001, 1003, 1005, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 8, 6, 16, 12, 22, 10, 38, 34, 14, 20, 58, 46, 26, 62, 18, 30, 52, 72, 102, 126, 24, 90, 68, 78, 28, 80, 138, 32, 150, 194, 84, 238, 36, 44, 94, 40, 220, 120, 42, 106, 88, 368, 250, 48, 288, 98, 50, 218, 208, 54, 432, 392, 56, 146, 160, 60, 324, 354, 188, 64, 268, 134, 66, 164, 156, 70, 244, 76, 184, 74, 360, 434, 436, 276, 236, 118, 278, 438, 82, 440, 142, 300, 86, 330, 442, 112, 444, 170, 92, 446, 262, 96, 352, 116, 166, 448, 100, 450, 132, 104, 212, 452, 322, 108, 388, 144, 110, 260, 206, 114, 256, 182, 454, 376, 294, 178, 350, 396, 122, 124, 298, 456, 200, 128, 316, 458, 130, 202, 340, -1, -1, 346, 136, 460, 176, 140, 462, 296, 234, -1, -1, 418, 464, 148, 466, -1, -1, 152, 468, 154, 230, 470, 344, 158, 304, 472, 198, 474, 162, -1, -1, 476, 306, 168, 478, -1, -1, 172, 480, 266, 174, -1, -1, 482, 484, 180, 332, -1, -1, -1, -1, 186, 366, -1, -1, 190, 486, 192, 488, -1, -1, 196, 356, 490, 492, -1, -1, 494, 496, 204, 498, -1, -1, -1, -1, 210, 500, -1, -1, 502, 214, 216, 504, -1, -1, 506, 508, 408, 222, 224, 334, 284, 226, 228, 510, 372, 308, 512, 232, -1, -1, -1, -1, -1, -1, 378, 240, 242, 364, 514, 342, 246, 338, 248, 362, -1, -1, 252, 516, 254, 518, -1, -1, 520, 258, -1, -1, -1, -1, 264, 522, -1, -1, -1, -1, 428, 270, 272, 310, 524, 274, 526, 528, -1, -1, 280, 404, 530, 282, -1, -1, 532, 286, 534, 536, 538, 290, 292, 414, 540, 370, -1, -1, -1, -1, 542, 544, 546, 302, -1, -1, 548, 550, 552, 554, -1, -1, 312, 556, 558, 314, -1, -1, 318, 560, 320, 562, 564, 566, 568, 570, 572, 326, 328, 574, 576, 578, -1, -1, -1, -1, 336, 580, 582, 584, 586, 588, 590, 592, 594, 596, -1, -1, 598, 348, 600, 374, 602, 604, 606, 608, 610, 612, 358, 614, -1, -1, 616, 618, -1, -1, 620, 622, -1, -1, 624, 626, -1, -1, -1, -1, -1, -1, -1, -1, 628, 380, 382, 384, 630, 632, 386, 634, -1, -1, 390, 636, 638, 640, 642, 394, 644, 646, 648, 398, 400, 650, 402, 652, -1, -1, 654, 406, -1, -1, 410, 420, 656, 412, 658, 660, 416, 662, -1, -1, -1, -1, 664, 422, 424, 666, 426, 668, -1, -1, 430, 670, 672, 674, 676, 678, 680, 682, 684, 686, 688, 690, -1, -1, -1, -1, 692, 694, 696, 698, 700, 702, -1, -1, 704, 706, -1, -1, 708, 710, 712, 714, 716, 718, 720, 722, -1, -1, -1, -1, 724, 726, -1, -1, -1, -1, -1, -1, 728, 730, -1, -1, 732, 734, -1, -1, -1, -1, 736, 738, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 740, 742, -1, -1, -1, -1, -1, -1, 744, 746, -1, -1, 748, 750, 752, 754, -1, -1, -1, -1, -1, -1, 756, 758, -1, -1, -1, -1, -1, -1, 760, 762, -1, -1, -1, -1, 764, 766, -1, -1, 768, 770, 772, 774, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 776, 778, -1, -1, 780, 782, 784, 786, -1, -1, -1, -1, -1, -1, -1, -1, 788, 790, 792, 794, -1, -1, -1, -1, 796, 798, 800, 802, 804, 806, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 808, 810, -1, -1, -1, -1, -1, -1, 812, 814, 816, 818, 820, 822, 824, 826, -1, -1, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 850, 852, 854, -1, -1, -1, -1, -1, -1, 856, 858, -1, -1, -1, -1, 860, 862, -1, -1, -1, -1, 864, 866, 868, 870, -1, -1, -1, -1, 872, 874, 876, 878, 880, 882, -1, -1, 884, 886, 888, 890, -1, -1, 892, 894, 896, 898, 900, 902, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, 952, 954, 956, 958, -1, -1, -1, -1, 960, 962, 964, 966, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, -1, -1, -1, -1, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, -1, -1, -1, -1, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 14, 18, 26, 10, 30, 40, 12, 44, 36, 50, 16, 78, 22, 20, 66, 62, 96, 24, 72, 60, 70, 28, 124, 142, 88, 32, 158, 114, 34, 232, 322, 180, 38, 58, 352, 418, 42, 48, 120, 46, 172, 92, 56, 224, 358, 52, 238, 152, 54, 84, 384, 166, 474, 268, 112, 138, 100, 64, 198, 476, 108, 192, 68, 202, 204, 86, 278, 186, 74, 76, 106, 228, 212, 80, 146, 118, 82, 478, 372, 378, 94, 480, 178, 262, 90, 382, 220, 308, 102, 104, 302, 482, 98, 282, 182, 156, 128, 136, 130, -1, -1, 314, 164, 484, 110, -1, -1, 214, 230, 462, 116, 270, 486, 134, 386, 122, 488, 252, 272, 290, 126, 132, 216, -1, -1, -1, -1, 490, 306, 492, 316, -1, -1, 376, 140, -1, -1, 334, 144, 494, 222, 148, 400, 496, 150, 250, 498, 424, 154, 500, 168, -1, -1, 160, 404, 340, 162, 328, 284, -1, -1, 208, 276, 374, 170, -1, -1, 428, 174, 394, 176, 502, 248, -1, -1, 504, 256, 184, 440, -1, -1, 366, 188, 190, 360, -1, -1, 194, 434, 370, 196, 266, 506, 508, 200, 380, 300, 346, 210, 296, 206, 510, 304, -1, -1, 512, 514, -1, -1, -1, -1, 218, 516, 390, 518, 520, 392, 522, 524, 362, 226, 526, 528, -1, -1, -1, -1, 530, 234, 236, 368, 532, 534, 444, 240, 242, 536, 458, 244, 538, 246, -1, -1, -1, -1, -1, -1, 254, 540, -1, -1, 258, 542, 398, 260, -1, -1, 264, 452, 544, 546, -1, -1, 350, 548, 550, 312, 274, 552, -1, -1, -1, -1, 280, 554, -1, -1, 556, 558, 286, 560, 288, 562, -1, -1, 292, 466, 318, 294, 564, 354, 298, 566, -1, -1, -1, -1, -1, -1, -1, -1, 568, 570, 310, 572, -1, -1, 574, 576, -1, -1, -1, -1, 578, 320, -1, -1, 324, 580, 326, 582, 584, 388, 586, 330, 332, 588, -1, -1, 590, 336, 338, 592, -1, -1, 594, 342, 344, 596, 356, 598, 348, 600, -1, -1, -1, -1, 602, 604, -1, -1, -1, -1, 606, 608, -1, -1, 364, 610, -1, -1, 612, 614, 416, 616, 618, 620, 622, 624, -1, -1, -1, -1, 456, 626, -1, -1, 628, 630, 632, 634, 636, 638, -1, -1, -1, -1, -1, -1, 396, 640, -1, -1, -1, -1, 402, 642, 644, 646, 406, 648, 650, 408, 410, 652, 414, 412, -1, -1, -1, -1, -1, -1, 654, 420, 422, 656, 658, 660, 662, 426, 664, 666, 668, 430, 442, 432, -1, -1, 436, 670, 672, 438, -1, -1, -1, -1, -1, -1, 470, 446, 674, 448, 450, 676, -1, -1, 678, 454, -1, -1, -1, -1, 460, 680, -1, -1, 682, 464, 684, 686, 688, 468, 690, 692, 694, 472, 696, 698, 700, 702, 704, 706, 708, 710, -1, -1, 712, 714, -1, -1, 716, 718, 720, 722, 724, 726, -1, -1, 728, 730, 732, 734, -1, -1, 736, 738, -1, -1, 740, 742, -1, -1, 744, 746, -1, -1, -1, -1, -1, -1, 748, 750, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 752, 754, -1, -1, -1, -1, 756, 758, -1, -1, -1, -1, 760, 762, -1, -1, -1, -1, -1, -1, 764, 766, -1, -1, -1, -1, -1, -1, -1, -1, 768, 770, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 772, 774, 776, 778, -1, -1, 780, 782, -1, -1, 784, 786, -1, -1, 788, 790, 792, 794, -1, -1, -1, -1, 796, 798, 800, 802, 804, 806, 808, 810, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 812, 814, 816, 818, -1, -1, -1, -1, -1, -1, 820, 822, -1, -1, -1, -1, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 850, 852, 854, -1, -1, -1, -1, 856, 858, 860, 862, -1, -1, 864, 866, -1, -1, -1, -1, -1, -1, 868, 870, 872, 874, 876, 878, 880, 882, -1, -1, -1, -1, 884, 886, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 888, 890, 892, 894, 896, 898, 900, 902, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 952, 954, 956, 958, 960, 962, 964, 966, -1, -1, -1, -1, 968, 970, 972, 974, 976, 978, 980, 982, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, 16, 18, 20, 22, 12, 14, 24, 26, 28, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90, 92, 94, 96, 98, 100, 102, 104, 106, 108, 110, 112, 114, 116, 118, 120, 122, 124, 126, 128, 130, 132, 134, 136, 138, 140, 142, 144, 146, 148, 150, 152, 154, 156, 158, 160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 180, 182, 184, 186, 188, 190, 192, 194, 196, 198, 200, 202, 204, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, 432, 434, 436, 438, 440, 442, 444, 446, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, 512, 514, 516, 518, 520, 522, 524, 526, 528, 530, 532, 534, 536, 538, 540, 542, 544, 546, 548, 550, 552, 554, 556, 558, 560, 562, 564, 566, 568, 570, 572, 574, 576, 578, 580, 582, 584, 586, 588, 590, 592, 594, 596, 598, 600, 602, 604, 606, 608, 610, 612, 614, 616, 618, 620, 622, 624, 626, 628, 630, 632, 634, 636, 638, 640, 642, 644, 646, 648, 650, 652, 654, 656, 658, 660, 662, 664, 666, 668, 670, 672, 674, 676, 678, 680, 682, 684, 686, 688, 690, 692, 694, 696, 698, 700, 702, 704, 706, 708, 710, 712, 714, 716, 718, 720, 722, 724, 726, 728, 730, 732, 734, 736, 738, 740, 742, 744, 746, 748, 750, 752, 754, 756, 758, 760, 762, 764, 766, 768, 770, 772, 774, 776, 778, 780, 782, 784, 786, 788, 790, 792, 794, 796, 798, 800, 802, 804, 806, 808, 810, 812, 814, 816, 818, 820, 822, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 850, 852, 854, 856, 858, 860, 862, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, 888, 890, 892, 894, 896, 898, 900, 902, 904, 906, 908, 910, 912, 914, 916, 918, 920, 922, 924, 926, 928, 930, 932, 934, 936, 938, 940, 942, 944, 946, 948, 950, 952, 954, 956, 958, 960, 962, 964, 966, 968, 970, 972, 974, 976, 978, 980, 982, 984, 986, 988, 990, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 5, 5, 10, 10, 4, 4, 16, 16, 11, 11, 6, 6, 22, 22, 14, 14, 26, 26, 17, 17, 29, 29, 9, 9, 34, 34, 8, 8, 37, 37, 40, 40, 35, 35, 13, 13, 45, 45, 48, 48, 18, 18, 51, 51, 54, 54, 12, 12, 57, 57, 15, 15, 61, 61, 64, 64, 24, 24, 67, 67, 19, 19, 71, 71, 69, 69, 25, 25, 27, 27, 80, 80, 32, 32, 84, 84, 42, 42, 23, 23, 90, 90, 36, 36, 93, 93, 47, 47, 98, 98, 20, 20, 101, 101, 41, 41, 105, 105, 108, 108, 87, 87, 111, 111, 95, 95, 77, 77, 39, 39, 120, 120, 121, 121, 21, 21, 125, 125, 128, 128, 100, 100, 63, 63, 134, 134, 28, 28, 137, 137, 82, 82, 107, 107, 55, 55, 145, 145, 30, 30, 149, 149, 151, 151, 66, 66, 155, 155, 56, 56, 160, 160, 65, 65, 96, 96, 165, 165, 89, 89, 169, 169, 172, 172, 136, 136, 117, 117, 177, 177, 113, 113, 70, 70, 183, 183, 60, 60, 187, 187, 189, 189, 31, 31, 193, 193, 158, 158, 124, 124, 129, 129, 201, 201, 110, 110, 50, 50, 207, 207, 102, 102, 212, 212, 213, 213, 49, 49, 38, 38, 220, 220, 221, 221, 224, 224, 225, 225, 152, 152, 230, 230, 140, 140, 76, 76, 33, 33, 238, 238, 239, 239, 68, 68, 243, 243, 245, 245, 44, 44, 249, 249, 251, 251, 112, 112, 256, 256, 109, 109, 92, 92, 261, 261, 171, 171, 62, 62, 268, 268, 269, 269, 272, 272, 75, 75, 78, 78, 277, 277, 280, 280, 223, 223, 284, 284, 46, 46, 288, 288, 289, 289, 116, 116, 139, 139, 122, 122, 83, 83, 300, 300, 156, 156, 164, 164, 228, 228, 270, 270, 309, 309, 312, 312, 126, 126, 315, 315, 317, 317, 104, 104, 58, 58, 324, 324, 325, 325, 85, 85, 178, 178, 222, 222, 333, 333, 244, 244, 130, 130, 242, 242, 154, 154, 133, 133, 346, 346, 118, 118, 94, 94, 59, 59, 194, 194, 355, 355, 72, 72, 246, 246, 240, 240, 184, 184, 43, 43, 292, 292, 227, 227, 348, 348, 115, 115, 237, 237, 378, 378, 379, 379, 380, 380, 383, 383, 106, 106, 387, 387, 53, 53, 392, 392, 119, 119, 396, 396, 397, 397, 399, 399, 278, 278, 404, 404, 219, 219, 407, 407, 410, 410, 290, 290, 413, 413, 143, 143, 408, 408, 420, 420, 421, 421, 423, 423, 267, 267, 427, 427, 52, 52, 73, 73, 74, 74, 79, 79, 81, 81, 86, 86, 88, 88, 91, 91, 97, 97, 99, 99, 103, 103, 114, 114, 123, 123, 127, 127, 135, 135, 138, 138, 144, 144, 146, 146, 150, 150, 153, 153, 157, 157, 159, 159, 163, 163, 166, 166, 170, 170, 175, 175, 176, 176, 188, 188, 190, 190, 195, 195, 196, 196, 199, 199, 200, 200, 202, 202, 208, 208, 211, 211, 214, 214, 217, 217, 218, 218, 226, 226, 229, 229, 241, 241, 250, 250, 252, 252, 255, 255, 262, 262, 271, 271, 273, 273, 274, 274, 279, 279, 283, 283, 285, 285, 286, 286, 287, 287, 291, 291, 297, 297, 298, 298, 299, 299, 303, 303, 304, 304, 305, 305, 306, 306, 310, 310, 311, 311, 316, 316, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 323, 323, 326, 326, 327, 327, 328, 328, 334, 334, 335, 335, 336, 336, 337, 337, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 345, 345, 347, 347, 349, 349, 350, 350, 351, 351, 352, 352, 353, 353, 354, 354, 356, 356, 359, 359, 360, 360, 363, 363, 364, 364, 367, 367, 368, 368, 377, 377, 381, 381, 382, 382, 384, 384, 388, 388, 389, 389, 390, 390, 391, 391, 393, 393, 394, 394, 395, 395, 398, 398, 400, 400, 403, 403, 409, 409, 411, 411, 412, 412, 414, 414, 419, 419, 422, 422, 424, 424, 428, 428, 429, 429, 430, 430, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 443, 443, 444, 444, 445, 445, 446, 446, 447, 447, 448, 448, 451, 451, 452, 452, 455, 455, 456, 456, 457, 457, 458, 458, 459, 459, 460, 460, 461, 461, 462, 462, 467, 467, 468, 468, 475, 475, 476, 476, 479, 479, 480, 480, 485, 485, 486, 486, 501, 501, 502, 502, 509, 509, 510, 510, 513, 513, 514, 514, 515, 515, 516, 516, 523, 523, 524, 524, 531, 531, 532, 532, 537, 537, 538, 538, 541, 541, 542, 542, 543, 543, 544, 544, 555, 555, 556, 556, 559, 559, 560, 560, 561, 561, 562, 562, 571, 571, 572, 572, 573, 573, 574, 574, 579, 579, 580, 580, 581, 581, 582, 582, 583, 583, 584, 584, 597, 597, 598, 598, 605, 605, 606, 606, 607, 607, 608, 608, 609, 609, 610, 610, 611, 611, 612, 612, 615, 615, 616, 616, 617, 617, 618, 618, 619, 619, 620, 620, 621, 621, 622, 622, 623, 623, 624, 624, 625, 625, 626, 626, 627, 627, 628, 628, 635, 635, 636, 636, 641, 641, 642, 642, 647, 647, 648, 648, 649, 649, 650, 650, 655, 655, 656, 656, 657, 657, 658, 658, 659, 659, 660, 660, 663, 663, 664, 664, 665, 665, 666, 666, 669, 669, 670, 670, 671, 671, 672, 672, 673, 673, 674, 674, 675, 675, 676, 676, 677, 677, 678, 678, 691, 691, 692, 692, 693, 693, 694, 694, 711, 711, 712, 712, 713, 713, 714, 714, 723, 723, 724, 724, 725, 725, 726, 726, 763, 763, 764, 764, 765, 765, 766, 766, 779, 779, 780, 780, 781, 781, 782, 782, 787, 787, 788, 788, 789, 789, 790, 790, 795, 795, 796, 796, 797, 797, 798, 798, 851, 851, 852, 852, 853, 853, 854, 854, 863, 863, 864, 864, 865, 865, 866, 866, 871, 871, 872, 872, 873, 873, 874, 874, 883, 883, 884, 884, 885, 885, 886, 886, 891, 891, 892, 892, 893, 893, 894, 894, 903, 903, 904, 904, 905, 905, 906, 906, 907, 907, 908, 908, 909, 909, 910, 910),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 10, 10, 4, 4, 14, 14, 5, 5, 17, 17, 16, 16, 21, 21, 6, 6, 25, 25, 8, 8, 29, 29, 32, 32, 12, 12, 36, 36, 9, 9, 40, 40, 11, 11, 43, 43, 41, 41, 13, 13, 49, 49, 52, 52, 46, 46, 37, 37, 23, 23, 19, 19, 61, 61, 18, 18, 66, 66, 24, 24, 22, 22, 72, 72, 73, 73, 15, 15, 77, 77, 80, 80, 53, 53, 69, 69, 28, 28, 88, 88, 45, 45, 84, 84, 20, 20, 96, 96, 60, 60, 92, 92, 93, 93, 74, 74, 64, 64, 108, 108, 58, 58, 31, 31, 114, 114, 79, 79, 42, 42, 119, 119, 26, 26, 124, 124, 100, 100, 102, 102, 125, 125, 117, 117, 101, 101, 59, 59, 138, 138, 27, 27, 142, 142, 78, 78, 145, 145, 148, 148, 51, 51, 152, 152, 99, 99, 30, 30, 157, 157, 160, 160, 106, 106, 55, 55, 154, 154, 168, 168, 44, 44, 172, 172, 174, 174, 86, 86, 35, 35, 98, 98, 181, 181, 71, 71, 186, 186, 187, 187, 65, 65, 191, 191, 194, 194, 62, 62, 198, 198, 67, 67, 68, 68, 204, 204, 165, 165, 202, 202, 76, 76, 111, 111, 126, 126, 215, 215, 90, 90, 144, 144, 47, 47, 224, 224, 75, 75, 112, 112, 33, 33, 232, 232, 233, 233, 50, 50, 238, 238, 239, 239, 242, 242, 244, 244, 176, 176, 149, 149, 121, 121, 251, 251, 180, 180, 255, 255, 258, 258, 87, 87, 261, 261, 195, 195, 57, 57, 115, 115, 122, 122, 271, 271, 166, 166, 70, 70, 277, 277, 97, 97, 162, 162, 283, 283, 285, 285, 123, 123, 289, 289, 292, 292, 203, 203, 295, 295, 200, 200, 94, 94, 206, 206, 132, 132, 91, 91, 307, 307, 270, 270, 105, 105, 134, 134, 291, 291, 318, 318, 34, 34, 321, 321, 323, 323, 161, 161, 328, 328, 329, 329, 141, 141, 334, 334, 335, 335, 159, 159, 340, 340, 341, 341, 201, 201, 345, 345, 267, 267, 38, 38, 294, 294, 343, 343, 48, 48, 188, 188, 223, 223, 361, 361, 185, 185, 234, 234, 193, 193, 82, 82, 167, 167, 137, 137, 83, 83, 199, 199, 89, 89, 54, 54, 118, 118, 326, 326, 217, 217, 220, 220, 173, 173, 393, 393, 257, 257, 146, 146, 399, 399, 158, 158, 403, 403, 406, 406, 407, 407, 410, 410, 409, 409, 367, 367, 39, 39, 418, 418, 419, 419, 151, 151, 424, 424, 171, 171, 428, 428, 430, 430, 192, 192, 433, 433, 436, 436, 182, 182, 429, 429, 237, 237, 444, 444, 446, 446, 447, 447, 262, 262, 452, 452, 377, 377, 241, 241, 457, 457, 113, 113, 462, 462, 290, 290, 466, 466, 443, 443, 470, 470, 56, 56, 63, 63, 81, 81, 85, 85, 95, 95, 107, 107, 116, 116, 120, 120, 131, 131, 133, 133, 143, 143, 147, 147, 150, 150, 153, 153, 175, 175, 179, 179, 196, 196, 197, 197, 205, 205, 209, 209, 210, 210, 216, 216, 218, 218, 219, 219, 221, 221, 222, 222, 225, 225, 226, 226, 231, 231, 235, 235, 236, 236, 240, 240, 243, 243, 252, 252, 256, 256, 263, 263, 264, 264, 268, 268, 269, 269, 272, 272, 278, 278, 281, 281, 282, 282, 284, 284, 286, 286, 293, 293, 296, 296, 305, 305, 306, 306, 308, 308, 311, 311, 312, 312, 317, 317, 322, 322, 324, 324, 325, 325, 327, 327, 330, 330, 333, 333, 336, 336, 339, 339, 342, 342, 344, 344, 346, 346, 351, 351, 352, 352, 357, 357, 358, 358, 362, 362, 365, 365, 366, 366, 368, 368, 369, 369, 370, 370, 371, 371, 372, 372, 378, 378, 381, 381, 382, 382, 383, 383, 384, 384, 385, 385, 386, 386, 394, 394, 400, 400, 401, 401, 402, 402, 404, 404, 405, 405, 408, 408, 417, 417, 420, 420, 421, 421, 422, 422, 423, 423, 425, 425, 426, 426, 427, 427, 434, 434, 435, 435, 445, 445, 448, 448, 451, 451, 458, 458, 461, 461, 463, 463, 464, 464, 465, 465, 467, 467, 468, 468, 469, 469, 471, 471, 472, 472, 473, 473, 474, 474, 475, 475, 476, 476, 477, 477, 478, 478, 481, 481, 482, 482, 485, 485, 486, 486, 487, 487, 488, 488, 489, 489, 490, 490, 493, 493, 494, 494, 495, 495, 496, 496, 499, 499, 500, 500, 503, 503, 504, 504, 507, 507, 508, 508, 515, 515, 516, 516, 529, 529, 530, 530, 535, 535, 536, 536, 541, 541, 542, 542, 549, 549, 550, 550, 559, 559, 560, 560, 579, 579, 580, 580, 581, 581, 582, 582, 585, 585, 586, 586, 589, 589, 590, 590, 593, 593, 594, 594, 595, 595, 596, 596, 601, 601, 602, 602, 603, 603, 604, 604, 605, 605, 606, 606, 607, 607, 608, 608, 631, 631, 632, 632, 633, 633, 634, 634, 641, 641, 642, 642, 647, 647, 648, 648, 649, 649, 650, 650, 651, 651, 652, 652, 653, 653, 654, 654, 655, 655, 656, 656, 657, 657, 658, 658, 659, 659, 660, 660, 661, 661, 662, 662, 667, 667, 668, 668, 669, 669, 670, 670, 673, 673, 674, 674, 681, 681, 682, 682, 683, 683, 684, 684, 685, 685, 686, 686, 687, 687, 688, 688, 693, 693, 694, 694, 711, 711, 712, 712, 713, 713, 714, 714, 715, 715, 716, 716, 717, 717, 718, 718, 719, 719, 720, 720, 721, 721, 722, 722, 739, 739, 740, 740, 741, 741, 742, 742, 751, 751, 752, 752, 753, 753, 754, 754, 755, 755, 756, 756, 757, 757, 758, 758, 771, 771, 772, 772, 773, 773, 774, 774, 787, 787, 788, 788, 789, 789, 790, 790, 823, 823, 824, 824, 825, 825, 826, 826, 827, 827, 828, 828, 829, 829, 830, 830, 835, 835, 836, 836, 837, 837, 838, 838, 839, 839, 840, 840, 841, 841, 842, 842, 867, 867, 868, 868, 869, 869, 870, 870, 951, 951, 952, 952, 953, 953, 954, 954, 955, 955, 956, 956, 957, 957, 958, 958, 967, 967, 968, 968, 969, 969, 970, 970, 971, 971, 972, 972, 973, 973, 974, 974),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10, 5, 5, 6, 6, 7, 7, 8, 8, 11, 11, 12, 12, 13, 13, 14, 14, 15, 15, 16, 16, 17, 17, 18, 18, 19, 19, 20, 20, 21, 21, 22, 22, 23, 23, 24, 24, 25, 25, 26, 26, 27, 27, 28, 28, 29, 29, 30, 30, 31, 31, 32, 32, 33, 33, 34, 34, 35, 35, 36, 36, 37, 37, 38, 38, 39, 39, 40, 40, 41, 41, 42, 42, 43, 43, 44, 44, 45, 45, 46, 46, 47, 47, 48, 48, 49, 49, 50, 50, 51, 51, 52, 52, 53, 53, 54, 54, 55, 55, 56, 56, 57, 57, 58, 58, 59, 59, 60, 60, 61, 61, 62, 62, 63, 63, 64, 64, 65, 65, 66, 66, 67, 67, 68, 68, 69, 69, 70, 70, 71, 71, 72, 72, 73, 73, 74, 74, 75, 75, 76, 76, 77, 77, 78, 78, 79, 79, 80, 80, 81, 81, 82, 82, 83, 83, 84, 84, 85, 85, 86, 86, 87, 87, 88, 88, 89, 89, 90, 90, 91, 91, 92, 92, 93, 93, 94, 94, 95, 95, 96, 96, 97, 97, 98, 98, 99, 99, 100, 100, 101, 101, 102, 102, 103, 103, 104, 104, 105, 105, 106, 106, 107, 107, 108, 108, 109, 109, 110, 110, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 117, 117, 118, 118, 119, 119, 120, 120, 121, 121, 122, 122, 123, 123, 124, 124, 125, 125, 126, 126, 127, 127, 128, 128, 129, 129, 130, 130, 131, 131, 132, 132, 133, 133, 134, 134, 135, 135, 136, 136, 137, 137, 138, 138, 139, 139, 140, 140, 141, 141, 142, 142, 143, 143, 144, 144, 145, 145, 146, 146, 147, 147, 148, 148, 149, 149, 150, 150, 151, 151, 152, 152, 153, 153, 154, 154, 155, 155, 156, 156, 157, 157, 158, 158, 159, 159, 160, 160, 161, 161, 162, 162, 163, 163, 164, 164, 165, 165, 166, 166, 167, 167, 168, 168, 169, 169, 170, 170, 171, 171, 172, 172, 173, 173, 174, 174, 175, 175, 176, 176, 177, 177, 178, 178, 179, 179, 180, 180, 181, 181, 182, 182, 183, 183, 184, 184, 185, 185, 186, 186, 187, 187, 188, 188, 189, 189, 190, 190, 191, 191, 192, 192, 193, 193, 194, 194, 195, 195, 196, 196, 197, 197, 198, 198, 199, 199, 200, 200, 201, 201, 202, 202, 203, 203, 204, 204, 205, 205, 206, 206, 207, 207, 208, 208, 209, 209, 210, 210, 211, 211, 212, 212, 213, 213, 214, 214, 215, 215, 216, 216, 217, 217, 218, 218, 219, 219, 220, 220, 221, 221, 222, 222, 223, 223, 224, 224, 225, 225, 226, 226, 227, 227, 228, 228, 229, 229, 230, 230, 231, 231, 232, 232, 233, 233, 234, 234, 235, 235, 236, 236, 237, 237, 238, 238, 239, 239, 240, 240, 241, 241, 242, 242, 243, 243, 244, 244, 245, 245, 246, 246, 247, 247, 248, 248, 249, 249, 250, 250, 251, 251, 252, 252, 253, 253, 254, 254, 255, 255, 256, 256, 257, 257, 258, 258, 259, 259, 260, 260, 261, 261, 262, 262, 263, 263, 264, 264, 265, 265, 266, 266, 267, 267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 272, 273, 273, 274, 274, 275, 275, 276, 276, 277, 277, 278, 278, 279, 279, 280, 280, 281, 281, 282, 282, 283, 283, 284, 284, 285, 285, 286, 286, 287, 287, 288, 288, 289, 289, 290, 290, 291, 291, 292, 292, 293, 293, 294, 294, 295, 295, 296, 296, 297, 297, 298, 298, 299, 299, 300, 300, 301, 301, 302, 302, 303, 303, 304, 304, 305, 305, 306, 306, 307, 307, 308, 308, 309, 309, 310, 310, 311, 311, 312, 312, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 323, 323, 324, 324, 325, 325, 326, 326, 327, 327, 328, 328, 329, 329, 330, 330, 331, 331, 332, 332, 333, 333, 334, 334, 335, 335, 336, 336, 337, 337, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 345, 345, 346, 346, 347, 347, 348, 348, 349, 349, 350, 350, 351, 351, 352, 352, 353, 353, 354, 354, 355, 355, 356, 356, 357, 357, 358, 358, 359, 359, 360, 360, 361, 361, 362, 362, 363, 363, 364, 364, 365, 365, 366, 366, 367, 367, 368, 368, 369, 369, 370, 370, 371, 371, 372, 372, 373, 373, 374, 374, 375, 375, 376, 376, 377, 377, 378, 378, 379, 379, 380, 380, 381, 381, 382, 382, 383, 383, 384, 384, 385, 385, 386, 386, 387, 387, 388, 388, 389, 389, 390, 390, 391, 391, 392, 392, 393, 393, 394, 394, 395, 395, 396, 396, 397, 397, 398, 398, 399, 399, 400, 400, 401, 401, 402, 402, 403, 403, 404, 404, 405, 405, 406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 412, 412, 413, 413, 414, 414, 415, 415, 416, 416, 417, 417, 418, 418, 419, 419, 420, 420, 421, 421, 422, 422, 423, 423, 424, 424, 425, 425, 426, 426, 427, 427, 428, 428, 429, 429, 430, 430, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446, 447, 447, 448, 448, 449, 449, 450, 450, 451, 451, 452, 452, 453, 453, 454, 454, 455, 455, 456, 456, 457, 457, 458, 458, 459, 459, 460, 460, 461, 461, 462, 462, 463, 463, 464, 464, 465, 465, 466, 466, 467, 467, 468, 468, 469, 469, 470, 470, 471, 471, 472, 472, 473, 473, 474, 474, 475, 475, 476, 476, 477, 477, 478, 478, 479, 479, 480, 480, 481, 481, 482, 482, 483, 483, 484, 484, 485, 485, 486, 486, 487, 487, 488, 488, 489, 489, 490, 490, 491, 491, 492, 492, 493, 493, 494, 494, 495, 495, 496, 496, 497, 497, 498, 498, 499, 499, 500, 500, 501, 501, 502, 502, 503, 503, 504, 504, 505, 505, 506, 506, 507, 507, 508, 508, 509, 509, 510, 510)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 3, 3, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 5, 5, 6, 6, 4, 4, 5, 5, 3, 3, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 7, 7, 5, 5, 6, 6, 7, 7, 5, 5, 6, 6, 4, 4, 5, 5, 6, 6, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 6, 6, 7, 7, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 7, 7, 5, 5, 6, 6, 7, 7, 5, 5, 6, 6, 7, 7, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 9, 9, 7, 7, 9, 9, 7, 7, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 6, 6, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 3, 3, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 4, 4, 5, 5, 3, 3, 4, 4, 5, 5, 5, 5, 6, 6, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 4, 4, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 6, 6, 7, 7, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 5, 5, 6, 6, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 9, 9, 4, 4, 5, 5, 6, 6, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 6, 6, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 7, 7, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 7, 7, 9, 9, 7, 7, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((131, 132, 141, 142, 147, 148, 161, 162, 167, 168, 173, 174, 179, 180, 181, 182, 185, 186, 191, 192, 197, 198, 203, 204, 205, 206, 209, 210, 215, 216, 231, 232, 233, 234, 235, 236, 247, 248, 253, 254, 257, 258, 259, 260, 263, 264, 265, 266, 275, 276, 281, 282, 293, 294, 295, 296, 301, 302, 307, 308, 313, 314, 329, 330, 331, 332, 343, 344, 357, 358, 361, 362, 365, 366, 369, 370, 371, 372, 373, 374, 375, 376, 385, 386, 401, 402, 405, 406, 415, 416, 417, 418, 425, 426, 439, 440, 441, 442, 449, 450, 453, 454, 463, 464, 465, 466, 469, 470, 471, 472, 473, 474, 477, 478, 481, 482, 483, 484, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 503, 504, 505, 506, 507, 508, 511, 512, 517, 518, 519, 520, 521, 522, 525, 526, 527, 528, 529, 530, 533, 534, 535, 536, 539, 540, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 557, 558, 563, 564, 565, 566, 567, 568, 569, 570, 575, 576, 577, 578, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 599, 600, 601, 602, 603, 604, 613, 614, 629, 630, 631, 632, 633, 634, 637, 638, 639, 640, 643, 644, 645, 646, 651, 652, 653, 654, 661, 662, 667, 668, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 715, 716, 717, 718, 719, 720, 721, 722, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 759, 760, 761, 762, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 783, 784, 785, 786, 791, 792, 793, 794, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 855, 856, 857, 858, 859, 860, 861, 862, 867, 868, 869, 870, 875, 876, 877, 878, 879, 880, 881, 882, 887, 888, 889, 890, 895, 896, 897, 898, 899, 900, 901, 902, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (103, 104, 109, 110, 127, 128, 129, 130, 135, 136, 139, 140, 155, 156, 163, 164, 169, 170, 177, 178, 183, 184, 189, 190, 207, 208, 211, 212, 213, 214, 227, 228, 229, 230, 245, 246, 247, 248, 249, 250, 253, 254, 259, 260, 265, 266, 273, 274, 275, 276, 279, 280, 287, 288, 297, 298, 299, 300, 301, 302, 303, 304, 309, 310, 313, 314, 315, 316, 319, 320, 331, 332, 337, 338, 347, 348, 349, 350, 353, 354, 355, 356, 359, 360, 363, 364, 373, 374, 375, 376, 379, 380, 387, 388, 389, 390, 391, 392, 395, 396, 397, 398, 411, 412, 413, 414, 415, 416, 431, 432, 437, 438, 439, 440, 441, 442, 449, 450, 453, 454, 455, 456, 459, 460, 479, 480, 483, 484, 491, 492, 497, 498, 501, 502, 505, 506, 509, 510, 511, 512, 513, 514, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 531, 532, 533, 534, 537, 538, 539, 540, 543, 544, 545, 546, 547, 548, 551, 552, 553, 554, 555, 556, 557, 558, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 583, 584, 587, 588, 591, 592, 597, 598, 599, 600, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 635, 636, 637, 638, 639, 640, 643, 644, 645, 646, 663, 664, 665, 666, 671, 672, 675, 676, 677, 678, 679, 680, 689, 690, 691, 692, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 723, 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 743, 744, 745, 746, 747, 748, 749, 750, 759, 760, 761, 762, 763, 764, 765, 766, 767, 768, 769, 770, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 831, 832, 833, 834, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 863, 864, 865, 866, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 959, 960, 961, 962, 963, 964, 965, 966, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 759, 760, 761, 762, 763, 764, 765, 766, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 863, 864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 1, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 2, 1, 1, 0, 1, 2, 1, 2, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 2, 0, 0, 2, 1, 1, 0, 2, 0, 1, 2, 0, 0, 0, 2, -2, 1, 1, 1, 0, -2, -2, -2, 1, 1, 1, 0, 0, 0, 2, 0, 1, 2, 2, 0, 0, 0, 1, 1, 0, -2, 0, 0, 2, 2, -2, 1, 0, 1, 2, -2, 1, 1, 1, 2, 0, 2, 1, 0, -2, 2, 0, -2, 2, -2, 1, 0, 1, 1, 1, 0, 1, 2, 1, -2, 0, 0, 0, 0, -2, 0, -2, 0, -2, -2, 1, 0, -2, 1, -2, -2, 1, 1, 2, 1, 1, -2, -2, -2, -2, 2, 1, 1, -2, -2, -2, -2, -2, 1, -2, -2, -2, 2, 0, 0, -2, -2, 1, 1, 0, -2, -2, -2, -2, -2, 1, 1, 1, 2, 1, 2, 1, -2, -2, 0, -2, -2, -2, -2, -2, 1, 1, -2, -2, -2, 1, 1, 2, 0, 1, 1, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, 2, 1, 1, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, -2, 0, 1, -2, -2, -2, -2, 1, -2, -2, -2, -2, 2, 0, 1, 0, 1, -2, -2, 0, -2, 2, 2, -2, 2, 0, 0, -2, -2, 1, 0, -2, -2, 0, -2, -2, -2, 1, 1, -2, 2, -2, -2, -2, -2, -2, 0, 1, -2, -2, -2, -2, 0, 0, -2, -2, -2, 0, -2, -2, 2, -2, -2, 0, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, 0, -2, 1, 0, -2, 1, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, 0, -2, 0, -2, -2, -2, 1, 0, 0, -2, -2, 2, -2, -2, 2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 0, 2, 0, 0, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, 1, -2, -2, -2, -2, 0, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, 0, -2, -2, -2, -2, 0, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 2, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 2, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, 2, 1, 2, 0, 2, 0, 0, 2, 2, 0, -2, 0, 0, 0, 0, -2, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, -2, 1, 0, 2, 1, 1, 1, 0, 1, 0, 2, 2, 1, -2, 1, 0, 1, 2, 2, 1, 0, 0, -2, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, -2, -2, 1, 1, -2, -2, 2, 0, 1, 1, 1, 2, 1, 0, -2, -2, 0, -2, 2, -2, -2, -2, 2, 1, 1, 2, -2, -2, 1, 0, 1, 0, -2, -2, -2, 0, -2, -2, 1, 2, 0, -2, 0, 1, 2, 2, 0, 1, -2, -2, 1, 0, 2, 0, -2, 0, 0, 0, 0, 1, 0, 2, 1, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, 0, -2, 0, -2, -2, 0, -2, -2, -2, 1, 1, 2, 1, 1, 0, -2, 1, 0, 0, -2, -2, -2, -2, 0, 0, -2, -2, -2, -2, 2, -2, 1, -2, -2, -2, -2, 1, -2, -2, -2, 2, -2, 1, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, 1, -2, 1, 2, -2, -2, 0, 0, -2, -2, -2, -2, -2, -2, 2, 1, -2, -2, 1, 0, -2, -2, 1, -2, -2, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, -2, 0, 1, 0, -2, -2, 1, -2, -2, -2, 1, -2, -2, 2, -2, 1, -2, -2, 0, -2, -2, -2, -2, 1, 0, 1, 2, 0, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 2, -2, 1, -2, -2, -2, 1, 1, 1, -2, -2, -2, -2, -2, -2, 2, -2, -2, -2, -2, -2, -2, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, 0, -2, 0, 2, -2, 0, -2, -2, 2, 1, -2, -2, -2, 2, 0, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 1, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, -2, 0, 2, -2, -2, -2, -2, 2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 0, -2, -2, 1, -2, -2, -2, -2, 1, -2, -2, 1, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, -2, -2, -2, -2, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((17096536, 894293, 27532130, 4500358, 11096038, 346653, 655327, 1354514, 35381898, 1201698, 68567, 1210534, 469637, 1458598, 1620590, 112505, 1882452, 9935275, 1164451, 56033, 1321223, 5230436, 7776885, 6689824, 9871128, 20862754, 21744058, 1014122, 68567, 1122188, 56033, 22807436, 19526907, 46858, 1297265, 1561604, 41955202, 1464762, 56033, 1721461, 68567, 1627674, 83804, 1446572, 1601748, 26331233, 1742961, 32282573, 1911925, 2686299, 4004811, 2633624, 46858, 13127936, 15107246, 68567, 1422893, 1170705, 13199456, 83804, 14777546, 919179, 46858, 23533789, 26814023, 21949093, 46858, -131072, 1442014, 1723956, 1794326, 325775, -131072, -131072, -131072, 212009, 288636, 176643, 1622828, 30147142, 31710530, 56033, 11255750, 777337, 68567, 83804, 18907520, 12646006, 11794382, 960731, 1068735, 12101702, -131072, 8557616, 9773811, 83804, 56033, -131072, 838379, 25049419, 1712166, 68567, -131072, 1515127, 1567105, 1388664, 46858, 33062855, 56033, 1526574, 34724178, -131072, 46858, 24270668, -131072, 46858, -131072, 1598362, 32149207, 1633735, 1619325, 525851, 5957636, 498430, 68567, 559337, -131072, 3162867, 3257396, 22296124, 18655202, -131072, 12982608, -131072, 14760109, -131072, -131072, 1211339, 15402974, -131072, 1282974, -131072, -131072, 1547983, 1555583, 56033, 1635929, 1497723, -131072, -131072, -131072, -131072, 56033, 1366672, 1415346, -131072, -131072, -131072, -131072, -131072, 1041045, -131072, -131072, -131072, 46858, 23380359, 23900357, -131072, -131072, 680748, 751089, 5188858, -131072, -131072, -131072, -131072, -131072, 1673518, 1792229, 1616435, 46858, 1718849, 56033, 1822267, -131072, -131072, 37365372, -131072, -131072, -131072, -131072, -131072, 388293, 1403152, -131072, -131072, -131072, 928387, 1043836, 68567, 10289857, 906891, 1003655, -131072, -131072, -131072, -131072, -131072, -131072, 943092, -131072, -131072, -131072, 68567, 1336365, 1319675, -131072, 1241434, -131072, -131072, -131072, -131072, 1227826, -131072, -131072, -131072, -131072, 3934948, 571078, -131072, -131072, -131072, -131072, 244720, -131072, -131072, -131072, -131072, 46858, 20626695, 1191680, 19344011, 1174759, -131072, -131072, 16325754, -131072, 83804, 68567, -131072, 83804, 21014326, 23048590, -131072, -131072, 798135, 7895337, -131072, -131072, 39244938, -131072, -131072, -131072, 819253, 859260, -131072, 56033, -131072, -131072, -131072, -131072, -131072, 33465809, 422876, -131072, -131072, -131072, -131072, 2284535, 2010488, -131072, -131072, -131072, 24240464, -131072, -131072, 56033, -131072, -131072, 16065858, -131072, -131072, -131072, -131072, -131072, 46858, -131072, -131072, -131072, -131072, 14325889, -131072, -131072, -131072, -131072, -131072, -131072, 2249523, -131072, 1563087, 36033382, -131072, 1619893, -131072, 37918266, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 24769735, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1082660, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 573678, -131072, -131072, 56033, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 46858, 29491787, -131072, 28842135, -131072, -131072, -131072, 926995, 9224948, 7992198, -131072, -131072, 56033, -131072, -131072, 83804, -131072, -131072, -131072, -131072, -131072, -131072, 427482, -131072, -131072, -131072, -131072, -131072, 45171106, 46858, 46151048, 44234234, -131072, -131072, -131072, 45860976, -131072, -131072, -131072, -131072, -131072, 677831, -131072, -131072, -131072, -131072, 1339435, -131072, -131072, 1157687, -131072, -131072, -131072, -131072, 3946753, -131072, -131072, 1592144, -131072, -131072, -131072, -131072, 1567361, -131072, -131072, -131072, 1192433, -131072, -131072, 29208879, -131072, -131072, -131072, -131072, 9237398, -131072, 974977, -131072, -131072, -131072, 861095, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072),
                (22349759, 839124, 32788236, 5769722, 15638489, 365977, 8050057, 1447213, 41229002, 1304261, 68567, 1563038, 1704790, 1073904, 1195395, 1058366, 68567, 1856382, 4544132, 133480, 2520230, 662456, 727899, 599323, 83804, 1286544, 1470781, 17533123, 21437198, 1196808, 46858, 30508610, 24304818, 22817571, 27852604, 83804, 28292616, 1631468, 44519502, 1547920, 56033, 46858, 34216624, 11611502, 13749468, 9756312, 56033, 881441, 68567, 15671868, 46858, 19992931, 17780119, 56033, 56033, 25492927, -131072, 29968826, 25710073, 341528, 1277260, -131072, 112986, 454420, 517990, 508949, 617281, 27545485, 24240684, 1468569, 1553952, 1674834, 37373628, 1672104, 1772762, 1315437, 18428466, 279921, 348351, -131072, 292001, 7876012, 68567, 919330, 984394, 974574, 11022837, 724085, 6839280, 46858, 46858, 1479627, -131072, 854829, 14019026, 1286185, 83804, 56033, 1336128, 20995669, 17168284, -131072, 19080953, 18053228, 1160082, 1579780, 29590895, 1632235, 1685640, 30563472, 32675447, 1563704, 1595924, 21617576, 1666028, 3116355, 4420363, 2502588, 46858, 928625, 999281, -131072, -131072, 1793187, 1895700, -131072, -131072, 56033, 26593368, 1396168, 1435144, 535393, 46858, 620894, 5961196, -131072, -131072, 7695402, -131072, 68567, -131072, -131072, -131072, 56033, 1181997, 1130144, 68567, -131072, -131072, 988404, 11863912, 960510, 12865776, -131072, -131072, -131072, 1011189, -131072, -131072, 1487106, 46858, 37244524, -131072, 35690168, 1618464, 68567, 83804, 5234918, 586795, -131072, -131072, 711290, 9343383, 46858, 11754012, -131072, 8608740, 38109430, 38856884, 34474668, 1747720, 3408006, 56033, 724094, -131072, -131072, 6229980, -131072, -131072, -131072, 1498998, -131072, -131072, -131072, 25035322, -131072, 20808420, -131072, -131072, 8476939, -131072, -131072, -131072, 1201410, 1241648, 68567, 1316943, 1133725, 13853212, -131072, 1336215, 26846270, 29504202, -131072, -131072, -131072, -131072, 19603286, 20474830, -131072, -131072, -131072, -131072, 46858, -131072, 799849, -131072, -131072, -131072, -131072, 1113159, -131072, -131072, -131072, 68567, -131072, 892906, -131072, -131072, 56033, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1642067, -131072, 1624466, 83804, -131072, -131072, 27154012, 28819401, -131072, -131072, -131072, -131072, -131072, -131072, 83804, 1421808, -131072, -131072, 1213760, 21676102, -131072, -131072, 1382145, -131072, -131072, -131072, -131072, -131072, 1459249, 26183500, -131072, -131072, -131072, -131072, -131072, -131072, 21656072, 1381228, 20767261, -131072, -131072, 1601150, -131072, -131072, -131072, 208349, -131072, -131072, 68567, -131072, 1775893, -131072, -131072, 33424657, -131072, -131072, -131072, -131072, 1733213, 45767622, 1724822, 46858, 43156564, -131072, -131072, -131072, -131072, -131072, -131072, 15783446, -131072, -131072, -131072, 1812901, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1718731, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 907675, -131072, -131072, -131072, -131072, -131072, 56033, -131072, 1352922, -131072, -131072, -131072, 510779, 583356, 546286, -131072, -131072, -131072, -131072, -131072, -131072, 56033, -131072, -131072, -131072, -131072, -131072, -131072, 38368630, 40739800, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1033587, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 40932084, -131072, -131072, -131072, 1725959, -131072, -131072, 12314512, -131072, 10401144, 68567, -131072, 13010510, -131072, -131072, 46858, 1046032, -131072, -131072, -131072, 46858, 6513634, -131072, -131072, -131072, -131072, 352310, -131072, -131072, -131072, -131072, -131072, 702083, -131072, -131072, -131072, 19278208, -131072, -131072, -131072, -131072, -131072, -131072, -131072, 1047452, -131072, -131072, -131072, -131072, 30760648, -131072, -131072, -131072, 508460, -131072, -131072, -131072, -131072, 23513862, 46858, -131072, -131072, -131072, -131072, 83804, -131072, -131072, -131072, -131072, 1309628, -131072, -131072, -131072, -131072, 9183654, -131072, -131072, 1380621, -131072, -131072, -131072, -131072, 1488939, -131072, -131072, 1818255, -131072, -131072, 1875076, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072),
                (33324485, 843327, 44551630, 8684409, 19000801, -131072, -131072, -131072, -131072, 1598180, 46202880, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072, -131072)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((19693, 9109, 21291, 16544, 1846, 6932, 20165, 17315, 21691, 21225, 6385, 14698, 1787, 1751, 13312, 3310, 19709, 199, 4912, 14461, 1430, 21588, 15964, 3236, 20144, 18072, 6927, 7412, 19051, 21754, 16908, 11776, 20913, 4228, 18866, 20286, 21807, 21650, 12726, 2764, 19136, 317, 11727, 11235, 21263, 5006, 18592, 13485, 21722, 6480, 294, 560, 18022, 13190, 2222, 5097, 328, 428, 11203, 2648, 17476, 4161, 19115, 6132, 665, 1820, 13523, 0, 20285, 9175, 20436, 9930, 0, 0, 21845, 14135, 21343, 21141, 3277, 14824, 1986, 16020, 21301, 8875, 19962, 17800, 7112, 14683, 21452, 6242, 19115, 18725, 0, 15420, 1456, 1298, 8995, 0, 16097, 1820, 14564, 20389, 0, 1214, 11360, 21806, 18826, 7282, 21625, 1365, 19115, 21845, 13653, 8738, 21845, 4681, 0, 496, 8091, 2819, 15197, 18893, 21787, 21605, 6554, 2731, 21845, 9709, 20436, 705, 7752, 16384, 1285, 21845, 12743, 0, 21845, 13107, 20972, 0, 10448, 14135, 0, 311, 4599, 11916, 1618, 6242, 21845, 15019, 4855, 0, 6242, 1456, 18204, 0, 13107, 10082, 18933, 0, 6242, 21845, 10194, 16384, 3855, 21092, 14564, 6242, 19859, 266, 5749, 13653, 0, 0, 21845, 21845, 9362, 21379, 21839, 21782, 17496, 1680, 20981, 17821, 21845, 21845, 10082, 0, 18725, 9362, 19661, 0, 14564, 14043, 21845, 17873, 0, 61, 1604, 10486, 144, 1820, 18485, 14564, 0, 21845, 12850, 10923, 0, 15124, 21845, 21845, 7282, 18303, 21673, 11763, 21845, 16991, 0, 21845, 7282, 0, 6242, 16384, 2185, 0, 6554, 63, 3799, 17476, 0, 6242, 0, 1365, 10923, 0, 8192, 21845, 20454, 14564, 21677, 4369, 20560, 0, 10923, 1755, 0, 705, 6899, 0, 18725, 21685, 17164, 8738, 21845, 16705, 21313, 20025, 8738, 5461, 0, 0, 13107, 19661, 21758, 21845, 14564, 6554, 21845, 21845, 13107, 21845, 15604, 15604, 21845, 21845, 7282, 21845, 19115, 7282, 21845, 14564, 0, 1702, 0, 0, 6242, 0, 16384, 4369, 0, 0, 10923, 21845, 13107, 5461, 0, 21845, 14564, 0, 2979, 0, 9362, 0, 7282, 0, 8738, 291, 7282, 21824, 20197, 7282, 20972, 14564, 21381, 0, 7282, 21845, 14564, 7282, 0, 7282, 0, 0, 7282, 7282, 0, 21845, 16384, 5461, 0, 20972, 14564, 21845, 16384, 21845, 14564, 1150, 7282, 21845, 14564, 14564, 21845, 0, 5461, 19418, 21845, 21845, 10923, 17476, 21845, 21845, 14564, 20954, 21845, 21845, 13107, 0, 21845, 4369, 0, 17476, 21845, 18204, 21845, 21845, 21141, 18204, 21845, 9362, 21845, 14564, 5461, 898, 25, 312, 14564, 0, 2731, 0, 7282, 19418, 21845, 14564, 21845, 18725, 21845, 0, 2427, 7282, 0, 19661, 21845, 21845, 21653, 17583, 21823, 2427, 21845, 0, 7282, 20025, 21845, 21845, 14564, 19418, 21845, 1820, 0, 0, 7282, 21845, 20165, 14564, 21845, 1560, 0, 7282, 0, 0, 1456, 7282, 0, 1820, 0, 0, 7282, 21845, 21221, 13107, 21845, 21845, 20632, 14564, 21845, 20632, 21845, 14564, 21845, 0, 364, 7282, 187, 5461, 0, 21845, 21203, 14564, 21845, 14564, 16384, 0, 0, 0, 0, 0, 0, 21845, 21845, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 16384, 16384, 21845, 21845, 0, 0, 21845, 21845, 0, 0, 0, 0, 16384, 16384, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 10923, 10923, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 17476, 17476, 0, 0, 10923, 10923, 21845, 21845, 0, 0, 10923, 10923, 0, 0, 0, 0, 8738, 8738, 21845, 21845, 0, 0, 0, 0, 13107, 13107, 21845, 21845, 21845, 21845, 13107, 13107, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 10923, 10923, 0, 0, 21845, 21845, 14564, 14564, 0, 0, 0, 0, 7282, 7282, 7282, 7282, 7282, 7282, 14564, 14564, 21845, 21845, 14564, 14564, 7282, 7282, 0, 0, 21845, 21845, 16384, 16384, 5461, 5461, 0, 0, 14564, 14564, 21845, 21845, 16384, 16384, 21845, 21845, 14564, 14564, 0, 0, 5461, 5461, 21845, 21845, 21845, 21845, 10923, 10923, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 0, 0, 0, 0, 7282, 7282, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 7282, 7282, 21845, 21845, 21845, 21845, 14564, 14564, 0, 0, 21845, 21845, 14564, 14564, 21845, 21845, 0, 0, 7282, 7282, 0, 0, 0, 0, 7282, 7282, 0, 0, 0, 0, 21845, 21845, 13107, 13107, 21845, 21845, 21845, 21845, 14564, 14564, 21845, 21845, 21845, 21845, 14564, 14564, 21845, 21845, 0, 0, 7282, 7282, 5461, 5461, 0, 0, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 17476, 17476, 17476, 17476, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 13107, 13107, 13107, 13107, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 16384, 16384, 16384, 16384, 5461, 5461, 5461, 5461, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 7282, 7282, 7282, 7282, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 7282, 7282, 7282, 7282, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845),
                (17504, 6471, 21131, 14934, 2088, 4995, 20596, 16572, 21686, 21205, 6171, 2265, 16575, 705, 6267, 18982, 2644, 11781, 1569, 3281, 20101, 15619, 21580, 20984, 3925, 662, 6522, 17417, 1794, 21817, 16634, 5534, 20238, 20747, 11083, 5273, 21400, 20196, 21828, 21682, 11792, 3624, 21373, 2752, 162, 822, 12629, 5521, 19034, 21587, 14794, 6117, 18811, 6117, 1060, 2427, 21845, 3641, 13544, 9029, 553, 0, 18811, 767, 6311, 21117, 2081, 767, 13835, 5461, 21005, 516, 8010, 2731, 16705, 11146, 20521, 13981, 21729, 21845, 1150, 277, 4896, 830, 13580, 20852, 2913, 2205, 13797, 1680, 10592, 4965, 21845, 17873, 3823, 20389, 7068, 4577, 179, 1150, 13559, 0, 18725, 2427, 15604, 49, 3396, 923, 10280, 19765, 3641, 910, 6595, 19859, 3121, 3750, 164, 408, 16991, 1150, 10448, 19661, 3361, 5461, 19418, 1214, 13653, 15391, 21378, 5461, 21065, 21672, 14564, 3121, 18569, 15604, 0, 6866, 0, 3766, 21845, 910, 17476, 15049, 21499, 7710, 19505, 18725, 0, 14947, 21499, 19859, 8192, 0, 16384, 21845, 9709, 0, 21845, 21835, 18858, 10923, 21845, 2570, 20389, 7282, 280, 3277, 18725, 5461, 21845, 21833, 20050, 10240, 21257, 0, 16384, 20753, 10923, 12483, 1337, 7282, 19765, 9102, 21845, 21845, 4855, 9102, 728, 16384, 3277, 3641, 16384, 7282, 20976, 21845, 9362, 21845, 7282, 11916, 21845, 21845, 6242, 50, 1090, 5345, 56, 1456, 20696, 0, 5461, 18204, 1986, 7282, 21845, 2427, 14564, 3121, 291, 892, 10923, 0, 10923, 18787, 21845, 10082, 21845, 18725, 0, 0, 6722, 17476, 0, 0, 1793, 0, 5861, 21845, 1986, 4749, 0, 0, 13653, 10923, 0, 0, 10923, 18725, 21845, 21239, 11763, 5461, 21845, 4201, 188, 0, 12136, 0, 8192, 0, 14564, 17476, 21550, 10923, 21845, 336, 5958, 10923, 0, 8738, 0, 3121, 21845, 15292, 21845, 331, 3427, 705, 7646, 14564, 21845, 0, 10923, 1900, 28, 683, 17476, 0, 7282, 4369, 0, 0, 2819, 17476, 0, 19275, 21845, 15604, 21845, 21845, 9362, 0, 4855, 15604, 21845, 21414, 21844, 21822, 15650, 2081, 21845, 5461, 446, 21845, 16384, 14564, 21671, 14564, 21845, 0, 5461, 10923, 0, 16384, 21845, 21845, 14564, 5461, 14564, 21845, 14564, 7282, 16384, 21845, 14564, 7282, 1560, 405, 7282, 7282, 0, 14564, 21845, 21845, 14564, 2731, 0, 1040, 14564, 0, 2185, 19986, 21845, 16991, 21845, 21845, 13902, 69, 1928, 8192, 0, 5461, 0, 21845, 16384, 0, 2570, 0, 5461, 0, 7282, 21845, 14564, 2731, 197, 0, 10923, 21845, 16384, 14564, 21845, 16384, 21845, 21845, 18204, 18725, 21845, 21845, 14564, 10923, 5461, 18204, 21845, 0, 2731, 7282, 0, 21845, 19418, 14564, 21845, 308, 0, 75, 2885, 0, 13902, 18725, 5461, 19418, 21755, 14564, 21845, 21845, 20665, 16384, 21845, 7282, 21845, 21845, 19859, 14564, 21845, 2185, 0, 0, 1820, 7282, 0, 21845, 20025, 14564, 21845, 1560, 0, 0, 1365, 21845, 20696, 14564, 21845, 7282, 10923, 1040, 0, 0, 7282, 539, 0, 280, 7282, 21845, 21504, 18569, 21845, 0, 21845, 0, 514, 0, 5461, 21845, 20696, 624, 0, 0, 7282, 21845, 21285, 14564, 21845, 326, 0, 0, 5461, 21845, 21554, 14564, 21845, 21731, 21845, 21845, 16384, 7282, 21845, 7282, 7282, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 5461, 5461, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 16384, 16384, 7282, 7282, 21845, 21845, 21845, 21845, 0, 0, 7282, 7282, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 0, 0, 17476, 17476, 0, 0, 0, 0, 17476, 17476, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 21845, 21845, 0, 0, 10923, 10923, 0, 0, 21845, 21845, 14564, 14564, 21845, 21845, 14564, 14564, 21845, 21845, 14564, 14564, 7282, 7282, 7282, 7282, 0, 0, 14564, 14564, 21845, 21845, 21845, 21845, 14564, 14564, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 7282, 7282, 0, 0, 10923, 10923, 21845, 21845, 0, 0, 21845, 21845, 14564, 14564, 21845, 21845, 0, 0, 0, 0, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 21845, 21845, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 7282, 7282, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 21845, 21845, 0, 0, 0, 0, 0, 0, 7282, 7282, 21845, 21845, 14564, 14564, 21845, 21845, 0, 0, 21845, 21845, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 7282, 7282, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 7282, 7282, 7282, 7282, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 7282, 7282, 7282, 7282, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 7282, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 14564, 14564, 14564, 14564, 14564, 14564, 14564, 14564, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 0, 0, 0, 0, 0, 0, 0, 0, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845),
                (10894, 3272, 21261, 9965, 1396, 2784, 21357, 355, 4823, 17674, 21835, 21653, 7341, 21294, 21845, 2784, 2784, 21357, 21357, 355, 355, 4823, 4823, 21653, 21653, 7341, 7341, 21294, 21294, 21845, 21845, 2784, 2784, 2784, 2784, 21357, 21357, 21357, 21357, 355, 355, 355, 355, 4823, 4823, 4823, 4823, 21653, 21653, 21653, 21653, 7341, 7341, 7341, 7341, 21294, 21294, 21294, 21294, 21845, 21845, 21845, 21845, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 355, 355, 355, 355, 355, 355, 355, 355, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 2784, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 21357, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 355, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 4823, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 21653, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 7341, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21294, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845, 21845)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 7, 5, 17, 11, 21, 9, 35, 29, 13, 15, 49, 63, 25, 71, 75, 197, 19, 27, 55, 121, 23, 95, 81, 43, 41, 53, 87, 237, 31, 33, 213, 129, 111, 37, 177, 105, 39, 115, 47, 329, 45, 85, 251, 99, 165, 69, 297, 51, 227, 307, 127, 61, 159, 57, 245, 289, 59, 221, 137, 131, 209, 65, 143, 151, 67, 451, 331, 79, 271, 73, 453, 455, 457, 77, 277, 333, 233, 157, 337, 83, 263, 93, 255, 193, 103, 89, 345, 91, 133, 339, 459, 189, 323, 169, 97, 461, 101, 225, 175, 361, 463, 359, 149, 365, 107, 109, 435, 343, 335, 465, 113, 155, 467, 117, 469, 423, 119, 231, 205, 123, 353, 327, 125, 207, 471, 191, 273, 303, 139, 473, 315, 475, 135, -1, -1, 161, 385, 477, 141, -1, -1, 283, 145, 147, 295, 203, 479, -1, -1, 481, 153, 321, 351, -1, -1, -1, -1, 483, 163, -1, -1, 485, 235, 405, 167, -1, -1, 407, 171, 173, 487, -1, -1, -1, -1, 179, 393, 309, 181, 259, 183, 185, 489, 491, 187, -1, -1, -1, -1, 493, 219, 195, 495, -1, -1, 373, 199, 201, 415, 325, 269, -1, -1, -1, -1, 497, 499, 211, 501, -1, -1, 215, 411, 217, 503, 293, 505, -1, -1, 507, 223, -1, -1, -1, -1, 419, 229, 509, 511, -1, -1, 319, 513, -1, -1, 515, 239, 241, 431, 243, 317, 517, 519, 247, 521, 299, 249, 523, 341, 381, 253, 525, 527, 257, 349, -1, -1, 261, 529, 531, 533, 265, 445, 535, 267, -1, -1, 537, 539, 541, 449, 275, 543, -1, -1, 545, 279, 281, 547, -1, -1, 285, 549, 551, 287, -1, -1, 291, 553, 555, 557, -1, -1, 305, 559, 561, 563, 565, 301, -1, -1, 567, 569, -1, -1, 387, 571, 427, 311, 573, 313, 575, 391, -1, -1, 577, 579, -1, -1, -1, -1, -1, -1, 581, 583, 585, 587, 589, 591, 363, 593, 595, 597, 599, 601, -1, -1, -1, -1, -1, -1, 603, 605, 347, 607, 609, 611, -1, -1, -1, -1, 355, 613, 615, 357, 617, 619, -1, -1, -1, -1, -1, -1, 621, 367, 369, 623, 371, 625, -1, -1, 375, 439, 377, 627, 629, 379, 631, 633, 383, 635, -1, -1, -1, -1, 637, 389, -1, -1, -1, -1, 639, 395, 397, 401, 399, 641, 643, 645, 403, 647, 649, 651, -1, -1, 409, 653, -1, -1, 655, 413, 657, 659, 417, 661, 663, 665, 667, 421, 669, 671, 425, 673, -1, -1, 675, 429, 677, 679, 681, 433, 683, 685, 437, 687, 689, 691, 693, 441, 695, 443, 697, 699, 701, 447, -1, -1, -1, -1, 703, 705, 707, 709, 711, 713, 715, 717, -1, -1, 719, 721, -1, -1, 723, 725, -1, -1, 727, 729, 731, 733, -1, -1, -1, -1, -1, -1, -1, -1, 735, 737, 739, 741, -1, -1, -1, -1, 743, 745, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 747, 749, -1, -1, -1, -1, 751, 753, 755, 757, -1, -1, 759, 761, -1, -1, -1, -1, 763, 765, -1, -1, -1, -1, -1, -1, 767, 769, -1, -1, -1, -1, -1, -1, 771, 773, 775, 777, -1, -1, -1, -1, 779, 781, -1, -1, 783, 785, -1, -1, 787, 789, -1, -1, -1, -1, -1, -1, 791, 793, 795, 797, -1, -1, -1, -1, -1, -1, 799, 801, 803, 805, -1, -1, -1, -1, -1, -1, 807, 809, 811, 813, 815, 817, 819, 821, 823, 825, 827, 829, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 831, 833, -1, -1, -1, -1, 835, 837, 839, 841, -1, -1, -1, -1, 843, 845, 847, 849, -1, -1, 851, 853, 855, 857, -1, -1, -1, -1, -1, -1, -1, -1, 859, 861, 863, 865, -1, -1, -1, -1, 867, 869, -1, -1, -1, -1, -1, -1, 871, 873, -1, -1, -1, -1, 875, 877, 879, 881, 883, 885, 887, 889, -1, -1, -1, -1, -1, -1, 891, 893, -1, -1, -1, -1, 895, 897, -1, -1, -1, -1, 899, 901, -1, -1, -1, -1, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, 951, 953, 955, 957, -1, -1, -1, -1, 959, 961, 963, 965, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 13, 17, 21, 9, 37, 29, 11, 53, 33, 43, 15, 49, 25, 19, 63, 59, 77, 23, 171, 131, 87, 97, 27, 75, 111, 451, 31, 55, 127, 193, 35, 67, 317, 39, 305, 159, 41, 71, 295, 45, 203, 81, 47, 93, 149, 315, 51, 103, 143, 57, 105, 209, 487, 89, 69, 61, 291, 489, 155, 115, 65, 325, 165, 337, 123, 189, 333, 373, 73, 179, 177, 95, 261, 79, 419, 491, 339, 233, 83, 345, 85, 363, 245, 137, 183, 275, 91, 135, 493, 213, 119, 377, 125, 99, 283, 265, 101, 495, 279, 229, 195, 443, 107, 253, 109, 303, 215, 217, 113, 381, 187, 117, 357, 365, 181, 311, 121, -1, -1, 243, 197, -1, -1, 129, 351, 269, 329, 413, 133, 369, 169, -1, -1, 139, 497, 141, 499, -1, -1, 145, 429, 147, 273, -1, -1, 151, 385, 313, 153, -1, -1, 501, 157, -1, -1, 475, 161, 163, 503, 287, 343, 167, 425, 257, 371, 505, 507, 467, 173, 175, 223, 509, 199, 391, 191, 331, 289, 259, 323, 185, 511, 513, 281, -1, -1, 515, 335, -1, -1, 517, 247, 519, 327, -1, -1, 201, 521, -1, -1, 401, 205, 207, 463, 239, 341, 523, 211, 379, 221, 525, 527, -1, -1, 219, 349, -1, -1, -1, -1, 225, 529, 227, 531, -1, -1, 533, 231, -1, -1, 535, 235, 537, 237, -1, -1, 241, 539, -1, -1, -1, -1, -1, -1, 249, 541, 383, 251, -1, -1, 255, 435, -1, -1, -1, -1, -1, -1, 263, 461, -1, -1, 433, 267, -1, -1, 271, 543, -1, -1, -1, -1, 423, 277, -1, -1, -1, -1, -1, -1, 285, 471, 301, 545, 547, 485, -1, -1, 549, 293, 551, 553, 297, 555, 299, 557, 559, 441, -1, -1, -1, -1, 307, 479, 397, 309, 319, 561, -1, -1, -1, -1, 563, 409, 565, 567, 569, 321, 571, 573, -1, -1, 575, 577, -1, -1, 579, 581, -1, -1, 583, 585, -1, -1, 361, 587, 589, 591, 593, 595, 597, 599, 347, 601, -1, -1, -1, -1, 353, 603, 355, 605, -1, -1, 447, 359, 389, 607, -1, -1, -1, -1, 609, 367, -1, -1, 611, 613, -1, -1, 375, 393, 615, 617, -1, -1, -1, -1, -1, -1, -1, -1, 387, 619, -1, -1, -1, -1, -1, -1, 621, 395, -1, -1, 623, 399, 625, 627, 403, 629, 457, 405, 631, 407, -1, -1, 411, 437, 633, 635, 637, 415, 417, 639, -1, -1, 641, 421, 643, 645, -1, -1, 647, 427, -1, -1, 649, 431, -1, -1, -1, -1, -1, -1, 651, 439, -1, -1, -1, -1, 445, 653, 655, 657, 449, 659, -1, -1, 661, 453, 455, 663, 665, 667, 669, 459, -1, -1, -1, -1, 465, 671, 673, 675, 677, 469, 679, 681, 473, 683, -1, -1, 685, 477, 687, 689, 481, 691, 693, 483, 695, 697, -1, -1, 699, 701, 703, 705, 707, 709, -1, -1, -1, -1, 711, 713, -1, -1, -1, -1, 715, 717, -1, -1, -1, -1, 719, 721, 723, 725, -1, -1, -1, -1, 727, 729, -1, -1, -1, -1, 731, 733, -1, -1, -1, -1, 735, 737, -1, -1, -1, -1, 739, 741, -1, -1, -1, -1, 743, 745, -1, -1, -1, -1, -1, -1, 747, 749, -1, -1, -1, -1, 751, 753, 755, 757, -1, -1, 759, 761, 763, 765, 767, 769, 771, 773, 775, 777, -1, -1, -1, -1, 779, 781, 783, 785, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 787, 789, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 791, 793, 795, 797, 799, 801, 803, 805, -1, -1, -1, -1, -1, -1, 807, 809, -1, -1, 811, 813, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 815, 817, -1, -1, -1, -1, -1, -1, 819, 821, 823, 825, 827, 829, 831, 833, -1, -1, 835, 837, -1, -1, -1, -1, 839, 841, 843, 845, 847, 849, -1, -1, 851, 853, 855, 857, 859, 861, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 887, 889, 891, 893, -1, -1, -1, -1, -1, -1, -1, -1, 895, 897, 899, 901, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 903, 905, 907, 909, -1, -1, -1, -1, 911, 913, 915, 917, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, 951, 953, 955, 957, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 959, 961, 963, 965, -1, -1, -1, -1, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, 15, 17, 19, 21, 11, 13, 23, 25, 27, 29, 31, 33, 35, 37, 39, 41, 43, 45, 47, 49, 51, 53, 55, 57, 59, 61, 63, 65, 67, 69, 71, 73, 75, 77, 79, 81, 83, 85, 87, 89, 91, 93, 95, 97, 99, 101, 103, 105, 107, 109, 111, 113, 115, 117, 119, 121, 123, 125, 127, 129, 131, 133, 135, 137, 139, 141, 143, 145, 147, 149, 151, 153, 155, 157, 159, 161, 163, 165, 167, 169, 171, 173, 175, 177, 179, 181, 183, 185, 187, 189, 191, 193, 195, 197, 199, 201, 203, 205, 207, 209, 211, 213, 215, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 237, 239, 241, 243, 245, 247, 249, 251, 253, 255, 257, 259, 261, 263, 265, 267, 269, 271, 273, 275, 277, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 341, 343, 345, 347, 349, 351, 353, 355, 357, 359, 361, 363, 365, 367, 369, 371, 373, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 415, 417, 419, 421, 423, 425, 427, 429, 431, 433, 435, 437, 439, 441, 443, 445, 447, 449, 451, 453, 455, 457, 459, 461, 463, 465, 467, 469, 471, 473, 475, 477, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, 511, 513, 515, 517, 519, 521, 523, 525, 527, 529, 531, 533, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 555, 557, 559, 561, 563, 565, 567, 569, 571, 573, 575, 577, 579, 581, 583, 585, 587, 589, 591, 593, 595, 597, 599, 601, 603, 605, 607, 609, 611, 613, 615, 617, 619, 621, 623, 625, 627, 629, 631, 633, 635, 637, 639, 641, 643, 645, 647, 649, 651, 653, 655, 657, 659, 661, 663, 665, 667, 669, 671, 673, 675, 677, 679, 681, 683, 685, 687, 689, 691, 693, 695, 697, 699, 701, 703, 705, 707, 709, 711, 713, 715, 717, 719, 721, 723, 725, 727, 729, 731, 733, 735, 737, 739, 741, 743, 745, 747, 749, 751, 753, 755, 757, 759, 761, 763, 765, 767, 769, 771, 773, 775, 777, 779, 781, 783, 785, 787, 789, 791, 793, 795, 797, 799, 801, 803, 805, 807, 809, 811, 813, 815, 817, 819, 821, 823, 825, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, 847, 849, 851, 853, 855, 857, 859, 861, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, 887, 889, 891, 893, 895, 897, 899, 901, 903, 905, 907, 909, 911, 913, 915, 917, 919, 921, 923, 925, 927, 929, 931, 933, 935, 937, 939, 941, 943, 945, 947, 949, 951, 953, 955, 957, 959, 961, 963, 965, 967, 969, 971, 973, 975, 977, 979, 981, 983, 985, 987, 989, 991, 993, 995, 997, 999, 1001, 1003, 1005, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 8, 6, 18, 12, 22, 10, 36, 30, 14, 16, 50, 64, 26, 72, 76, 198, 20, 28, 56, 122, 24, 96, 82, 44, 42, 54, 88, 238, 32, 34, 214, 130, 112, 38, 178, 106, 40, 116, 48, 330, 46, 86, 252, 100, 166, 70, 298, 52, 228, 308, 128, 62, 160, 58, 246, 290, 60, 222, 138, 132, 210, 66, 144, 152, 68, 452, 332, 80, 272, 74, 454, 456, 458, 78, 278, 334, 234, 158, 338, 84, 264, 94, 256, 194, 104, 90, 346, 92, 134, 340, 460, 190, 324, 170, 98, 462, 102, 226, 176, 362, 464, 360, 150, 366, 108, 110, 436, 344, 336, 466, 114, 156, 468, 118, 470, 424, 120, 232, 206, 124, 354, 328, 126, 208, 472, 192, 274, 304, 140, 474, 316, 476, 136, -1, -1, 162, 386, 478, 142, -1, -1, 284, 146, 148, 296, 204, 480, -1, -1, 482, 154, 322, 352, -1, -1, -1, -1, 484, 164, -1, -1, 486, 236, 406, 168, -1, -1, 408, 172, 174, 488, -1, -1, -1, -1, 180, 394, 310, 182, 260, 184, 186, 490, 492, 188, -1, -1, -1, -1, 494, 220, 196, 496, -1, -1, 374, 200, 202, 416, 326, 270, -1, -1, -1, -1, 498, 500, 212, 502, -1, -1, 216, 412, 218, 504, 294, 506, -1, -1, 508, 224, -1, -1, -1, -1, 420, 230, 510, 512, -1, -1, 320, 514, -1, -1, 516, 240, 242, 432, 244, 318, 518, 520, 248, 522, 300, 250, 524, 342, 382, 254, 526, 528, 258, 350, -1, -1, 262, 530, 532, 534, 266, 446, 536, 268, -1, -1, 538, 540, 542, 450, 276, 544, -1, -1, 546, 280, 282, 548, -1, -1, 286, 550, 552, 288, -1, -1, 292, 554, 556, 558, -1, -1, 306, 560, 562, 564, 566, 302, -1, -1, 568, 570, -1, -1, 388, 572, 428, 312, 574, 314, 576, 392, -1, -1, 578, 580, -1, -1, -1, -1, -1, -1, 582, 584, 586, 588, 590, 592, 364, 594, 596, 598, 600, 602, -1, -1, -1, -1, -1, -1, 604, 606, 348, 608, 610, 612, -1, -1, -1, -1, 356, 614, 616, 358, 618, 620, -1, -1, -1, -1, -1, -1, 622, 368, 370, 624, 372, 626, -1, -1, 376, 440, 378, 628, 630, 380, 632, 634, 384, 636, -1, -1, -1, -1, 638, 390, -1, -1, -1, -1, 640, 396, 398, 402, 400, 642, 644, 646, 404, 648, 650, 652, -1, -1, 410, 654, -1, -1, 656, 414, 658, 660, 418, 662, 664, 666, 668, 422, 670, 672, 426, 674, -1, -1, 676, 430, 678, 680, 682, 434, 684, 686, 438, 688, 690, 692, 694, 442, 696, 444, 698, 700, 702, 448, -1, -1, -1, -1, 704, 706, 708, 710, 712, 714, 716, 718, -1, -1, 720, 722, -1, -1, 724, 726, -1, -1, 728, 730, 732, 734, -1, -1, -1, -1, -1, -1, -1, -1, 736, 738, 740, 742, -1, -1, -1, -1, 744, 746, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 748, 750, -1, -1, -1, -1, 752, 754, 756, 758, -1, -1, 760, 762, -1, -1, -1, -1, 764, 766, -1, -1, -1, -1, -1, -1, 768, 770, -1, -1, -1, -1, -1, -1, 772, 774, 776, 778, -1, -1, -1, -1, 780, 782, -1, -1, 784, 786, -1, -1, 788, 790, -1, -1, -1, -1, -1, -1, 792, 794, 796, 798, -1, -1, -1, -1, -1, -1, 800, 802, 804, 806, -1, -1, -1, -1, -1, -1, 808, 810, 812, 814, 816, 818, 820, 822, 824, 826, 828, 830, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 832, 834, -1, -1, -1, -1, 836, 838, 840, 842, -1, -1, -1, -1, 844, 846, 848, 850, -1, -1, 852, 854, 856, 858, -1, -1, -1, -1, -1, -1, -1, -1, 860, 862, 864, 866, -1, -1, -1, -1, 868, 870, -1, -1, -1, -1, -1, -1, 872, 874, -1, -1, -1, -1, 876, 878, 880, 882, 884, 886, 888, 890, -1, -1, -1, -1, -1, -1, 892, 894, -1, -1, -1, -1, 896, 898, -1, -1, -1, -1, 900, 902, -1, -1, -1, -1, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, 952, 954, 956, 958, -1, -1, -1, -1, 960, 962, 964, 966, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 14, 18, 22, 10, 38, 30, 12, 54, 34, 44, 16, 50, 26, 20, 64, 60, 78, 24, 172, 132, 88, 98, 28, 76, 112, 452, 32, 56, 128, 194, 36, 68, 318, 40, 306, 160, 42, 72, 296, 46, 204, 82, 48, 94, 150, 316, 52, 104, 144, 58, 106, 210, 488, 90, 70, 62, 292, 490, 156, 116, 66, 326, 166, 338, 124, 190, 334, 374, 74, 180, 178, 96, 262, 80, 420, 492, 340, 234, 84, 346, 86, 364, 246, 138, 184, 276, 92, 136, 494, 214, 120, 378, 126, 100, 284, 266, 102, 496, 280, 230, 196, 444, 108, 254, 110, 304, 216, 218, 114, 382, 188, 118, 358, 366, 182, 312, 122, -1, -1, 244, 198, -1, -1, 130, 352, 270, 330, 414, 134, 370, 170, -1, -1, 140, 498, 142, 500, -1, -1, 146, 430, 148, 274, -1, -1, 152, 386, 314, 154, -1, -1, 502, 158, -1, -1, 476, 162, 164, 504, 288, 344, 168, 426, 258, 372, 506, 508, 468, 174, 176, 224, 510, 200, 392, 192, 332, 290, 260, 324, 186, 512, 514, 282, -1, -1, 516, 336, -1, -1, 518, 248, 520, 328, -1, -1, 202, 522, -1, -1, 402, 206, 208, 464, 240, 342, 524, 212, 380, 222, 526, 528, -1, -1, 220, 350, -1, -1, -1, -1, 226, 530, 228, 532, -1, -1, 534, 232, -1, -1, 536, 236, 538, 238, -1, -1, 242, 540, -1, -1, -1, -1, -1, -1, 250, 542, 384, 252, -1, -1, 256, 436, -1, -1, -1, -1, -1, -1, 264, 462, -1, -1, 434, 268, -1, -1, 272, 544, -1, -1, -1, -1, 424, 278, -1, -1, -1, -1, -1, -1, 286, 472, 302, 546, 548, 486, -1, -1, 550, 294, 552, 554, 298, 556, 300, 558, 560, 442, -1, -1, -1, -1, 308, 480, 398, 310, 320, 562, -1, -1, -1, -1, 564, 410, 566, 568, 570, 322, 572, 574, -1, -1, 576, 578, -1, -1, 580, 582, -1, -1, 584, 586, -1, -1, 362, 588, 590, 592, 594, 596, 598, 600, 348, 602, -1, -1, -1, -1, 354, 604, 356, 606, -1, -1, 448, 360, 390, 608, -1, -1, -1, -1, 610, 368, -1, -1, 612, 614, -1, -1, 376, 394, 616, 618, -1, -1, -1, -1, -1, -1, -1, -1, 388, 620, -1, -1, -1, -1, -1, -1, 622, 396, -1, -1, 624, 400, 626, 628, 404, 630, 458, 406, 632, 408, -1, -1, 412, 438, 634, 636, 638, 416, 418, 640, -1, -1, 642, 422, 644, 646, -1, -1, 648, 428, -1, -1, 650, 432, -1, -1, -1, -1, -1, -1, 652, 440, -1, -1, -1, -1, 446, 654, 656, 658, 450, 660, -1, -1, 662, 454, 456, 664, 666, 668, 670, 460, -1, -1, -1, -1, 466, 672, 674, 676, 678, 470, 680, 682, 474, 684, -1, -1, 686, 478, 688, 690, 482, 692, 694, 484, 696, 698, -1, -1, 700, 702, 704, 706, 708, 710, -1, -1, -1, -1, 712, 714, -1, -1, -1, -1, 716, 718, -1, -1, -1, -1, 720, 722, 724, 726, -1, -1, -1, -1, 728, 730, -1, -1, -1, -1, 732, 734, -1, -1, -1, -1, 736, 738, -1, -1, -1, -1, 740, 742, -1, -1, -1, -1, 744, 746, -1, -1, -1, -1, -1, -1, 748, 750, -1, -1, -1, -1, 752, 754, 756, 758, -1, -1, 760, 762, 764, 766, 768, 770, 772, 774, 776, 778, -1, -1, -1, -1, 780, 782, 784, 786, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 788, 790, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 792, 794, 796, 798, 800, 802, 804, 806, -1, -1, -1, -1, -1, -1, 808, 810, -1, -1, 812, 814, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 816, 818, -1, -1, -1, -1, -1, -1, 820, 822, 824, 826, 828, 830, 832, 834, -1, -1, 836, 838, -1, -1, -1, -1, 840, 842, 844, 846, 848, 850, -1, -1, 852, 854, 856, 858, 860, 862, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 888, 890, 892, 894, -1, -1, -1, -1, -1, -1, -1, -1, 896, 898, 900, 902, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 904, 906, 908, 910, -1, -1, -1, -1, 912, 914, 916, 918, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, 952, 954, 956, 958, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 960, 962, 964, 966, -1, -1, -1, -1, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, 16, 18, 20, 22, 12, 14, 24, 26, 28, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90, 92, 94, 96, 98, 100, 102, 104, 106, 108, 110, 112, 114, 116, 118, 120, 122, 124, 126, 128, 130, 132, 134, 136, 138, 140, 142, 144, 146, 148, 150, 152, 154, 156, 158, 160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 180, 182, 184, 186, 188, 190, 192, 194, 196, 198, 200, 202, 204, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, 432, 434, 436, 438, 440, 442, 444, 446, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, 512, 514, 516, 518, 520, 522, 524, 526, 528, 530, 532, 534, 536, 538, 540, 542, 544, 546, 548, 550, 552, 554, 556, 558, 560, 562, 564, 566, 568, 570, 572, 574, 576, 578, 580, 582, 584, 586, 588, 590, 592, 594, 596, 598, 600, 602, 604, 606, 608, 610, 612, 614, 616, 618, 620, 622, 624, 626, 628, 630, 632, 634, 636, 638, 640, 642, 644, 646, 648, 650, 652, 654, 656, 658, 660, 662, 664, 666, 668, 670, 672, 674, 676, 678, 680, 682, 684, 686, 688, 690, 692, 694, 696, 698, 700, 702, 704, 706, 708, 710, 712, 714, 716, 718, 720, 722, 724, 726, 728, 730, 732, 734, 736, 738, 740, 742, 744, 746, 748, 750, 752, 754, 756, 758, 760, 762, 764, 766, 768, 770, 772, 774, 776, 778, 780, 782, 784, 786, 788, 790, 792, 794, 796, 798, 800, 802, 804, 806, 808, 810, 812, 814, 816, 818, 820, 822, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 850, 852, 854, 856, 858, 860, 862, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, 888, 890, 892, 894, 896, 898, 900, 902, 904, 906, 908, 910, 912, 914, 916, 918, 920, 922, 924, 926, 928, 930, 932, 934, 936, 938, 940, 942, 944, 946, 948, 950, 952, 954, 956, 958, 960, 962, 964, 966, 968, 970, 972, 974, 976, 978, 980, 982, 984, 986, 988, 990, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 5, 5, 10, 10, 11, 11, 4, 4, 18, 18, 6, 6, 22, 22, 14, 14, 19, 19, 9, 9, 30, 30, 31, 31, 8, 8, 35, 35, 38, 38, 26, 26, 25, 25, 42, 42, 40, 40, 12, 12, 49, 49, 27, 27, 20, 20, 55, 55, 58, 58, 53, 53, 13, 13, 63, 63, 66, 66, 47, 47, 15, 15, 71, 71, 16, 16, 75, 75, 69, 69, 24, 24, 81, 81, 43, 43, 28, 28, 87, 87, 89, 89, 83, 83, 23, 23, 96, 96, 45, 45, 98, 98, 86, 86, 37, 37, 106, 106, 107, 107, 34, 34, 112, 112, 39, 39, 115, 115, 118, 118, 21, 21, 121, 121, 124, 124, 52, 52, 33, 33, 61, 61, 90, 90, 134, 134, 60, 60, 130, 130, 140, 140, 64, 64, 144, 144, 145, 145, 104, 104, 65, 65, 152, 152, 113, 113, 79, 79, 54, 54, 137, 137, 160, 160, 46, 46, 166, 166, 95, 95, 170, 170, 171, 171, 100, 100, 36, 36, 177, 177, 180, 180, 182, 182, 183, 183, 186, 186, 93, 93, 127, 127, 85, 85, 193, 193, 17, 17, 198, 198, 199, 199, 147, 147, 120, 120, 125, 125, 62, 62, 209, 209, 32, 32, 213, 213, 215, 215, 192, 192, 59, 59, 222, 222, 99, 99, 50, 50, 228, 228, 119, 119, 78, 78, 164, 164, 29, 29, 238, 238, 239, 239, 241, 241, 56, 56, 245, 245, 248, 248, 44, 44, 252, 252, 84, 84, 255, 255, 181, 181, 259, 259, 82, 82, 263, 263, 266, 266, 202, 202, 70, 70, 128, 128, 273, 273, 76, 76, 278, 278, 279, 279, 143, 143, 283, 283, 286, 286, 57, 57, 289, 289, 217, 217, 146, 146, 48, 48, 247, 247, 300, 300, 129, 129, 295, 295, 51, 51, 179, 179, 310, 310, 312, 312, 132, 132, 242, 242, 233, 233, 153, 153, 94, 94, 201, 201, 123, 123, 41, 41, 68, 68, 77, 77, 110, 110, 80, 80, 91, 91, 250, 250, 109, 109, 88, 88, 345, 345, 256, 256, 154, 154, 122, 122, 353, 353, 356, 356, 103, 103, 101, 101, 331, 331, 105, 105, 366, 366, 367, 367, 369, 369, 197, 197, 373, 373, 375, 375, 378, 378, 251, 251, 381, 381, 138, 138, 307, 307, 388, 388, 314, 314, 178, 178, 394, 394, 395, 395, 397, 397, 396, 396, 401, 401, 165, 165, 169, 169, 407, 407, 214, 214, 412, 412, 200, 200, 415, 415, 227, 227, 420, 420, 117, 117, 423, 423, 309, 309, 428, 428, 240, 240, 432, 432, 108, 108, 435, 435, 374, 374, 440, 440, 442, 442, 264, 264, 446, 446, 272, 272, 67, 67, 72, 72, 73, 73, 74, 74, 92, 92, 97, 97, 102, 102, 111, 111, 114, 114, 116, 116, 126, 126, 131, 131, 133, 133, 139, 139, 148, 148, 151, 151, 159, 159, 163, 163, 172, 172, 184, 184, 185, 185, 191, 191, 194, 194, 207, 207, 208, 208, 210, 210, 216, 216, 218, 218, 221, 221, 229, 229, 230, 230, 234, 234, 237, 237, 243, 243, 244, 244, 246, 246, 249, 249, 253, 253, 254, 254, 260, 260, 261, 261, 262, 262, 265, 265, 269, 269, 270, 270, 271, 271, 274, 274, 277, 277, 280, 280, 284, 284, 285, 285, 290, 290, 291, 291, 292, 292, 296, 296, 297, 297, 298, 298, 299, 299, 303, 303, 304, 304, 308, 308, 311, 311, 313, 313, 317, 317, 318, 318, 325, 325, 326, 326, 327, 327, 328, 328, 329, 329, 330, 330, 332, 332, 333, 333, 334, 334, 335, 335, 336, 336, 343, 343, 344, 344, 346, 346, 347, 347, 348, 348, 354, 354, 355, 355, 357, 357, 358, 358, 365, 365, 368, 368, 370, 370, 376, 376, 377, 377, 379, 379, 380, 380, 382, 382, 387, 387, 393, 393, 398, 398, 399, 399, 400, 400, 402, 402, 403, 403, 404, 404, 408, 408, 411, 411, 413, 413, 414, 414, 416, 416, 417, 417, 418, 418, 419, 419, 421, 421, 422, 422, 424, 424, 427, 427, 429, 429, 430, 430, 431, 431, 433, 433, 434, 434, 436, 436, 437, 437, 438, 438, 439, 439, 441, 441, 443, 443, 444, 444, 445, 445, 451, 451, 452, 452, 453, 453, 454, 454, 455, 455, 456, 456, 457, 457, 458, 458, 461, 461, 462, 462, 465, 465, 466, 466, 469, 469, 470, 470, 471, 471, 472, 472, 481, 481, 482, 482, 483, 483, 484, 484, 489, 489, 490, 490, 503, 503, 504, 504, 509, 509, 510, 510, 511, 511, 512, 512, 515, 515, 516, 516, 521, 521, 522, 522, 529, 529, 530, 530, 537, 537, 538, 538, 539, 539, 540, 540, 545, 545, 546, 546, 549, 549, 550, 550, 553, 553, 554, 554, 561, 561, 562, 562, 563, 563, 564, 564, 571, 571, 572, 572, 573, 573, 574, 574, 581, 581, 582, 582, 583, 583, 584, 584, 585, 585, 586, 586, 587, 587, 588, 588, 589, 589, 590, 590, 591, 591, 592, 592, 607, 607, 608, 608, 613, 613, 614, 614, 615, 615, 616, 616, 621, 621, 622, 622, 623, 623, 624, 624, 627, 627, 628, 628, 629, 629, 630, 630, 639, 639, 640, 640, 641, 641, 642, 642, 647, 647, 648, 648, 655, 655, 656, 656, 661, 661, 662, 662, 663, 663, 664, 664, 665, 665, 666, 666, 667, 667, 668, 668, 675, 675, 676, 676, 681, 681, 682, 682, 687, 687, 688, 688, 693, 693, 694, 694, 695, 695, 696, 696, 707, 707, 708, 708, 709, 709, 710, 710, 727, 727, 728, 728, 729, 729, 730, 730, 759, 759, 760, 760, 761, 761, 762, 762, 763, 763, 764, 764, 765, 765, 766, 766, 835, 835, 836, 836, 837, 837, 838, 838, 843, 843, 844, 844, 845, 845, 846, 846, 851, 851, 852, 852, 853, 853, 854, 854, 859, 859, 860, 860, 861, 861, 862, 862, 875, 875, 876, 876, 877, 877, 878, 878, 903, 903, 904, 904, 905, 905, 906, 906, 927, 927, 928, 928, 929, 929, 930, 930, 931, 931, 932, 932, 933, 933, 934, 934, 967, 967, 968, 968, 969, 969, 970, 970, 971, 971, 972, 972, 973, 973, 974, 974),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 10, 10, 4, 4, 14, 14, 5, 5, 17, 17, 6, 6, 21, 21, 16, 16, 26, 26, 9, 9, 30, 30, 12, 12, 34, 34, 8, 8, 37, 37, 40, 40, 13, 13, 43, 43, 46, 46, 15, 15, 50, 50, 11, 11, 31, 31, 53, 53, 19, 19, 59, 59, 18, 18, 64, 64, 35, 35, 58, 58, 41, 41, 72, 72, 27, 27, 20, 20, 77, 77, 45, 45, 82, 82, 84, 84, 24, 24, 57, 57, 90, 90, 47, 47, 75, 75, 25, 25, 97, 97, 100, 100, 51, 51, 54, 54, 106, 106, 108, 108, 28, 28, 112, 112, 63, 63, 115, 115, 94, 94, 120, 120, 68, 68, 96, 96, 32, 32, 127, 127, 23, 23, 132, 132, 91, 91, 87, 87, 137, 137, 139, 139, 52, 52, 143, 143, 145, 145, 48, 48, 149, 149, 152, 152, 62, 62, 156, 156, 39, 39, 160, 160, 161, 161, 66, 66, 165, 165, 134, 134, 22, 22, 172, 172, 173, 173, 74, 74, 73, 73, 118, 118, 88, 88, 183, 183, 114, 114, 69, 69, 178, 178, 33, 33, 104, 104, 124, 124, 176, 176, 199, 199, 44, 44, 204, 204, 205, 205, 55, 55, 210, 210, 93, 93, 110, 110, 111, 111, 217, 217, 212, 212, 174, 174, 223, 223, 225, 225, 103, 103, 230, 230, 81, 81, 234, 234, 236, 236, 207, 207, 239, 239, 123, 123, 86, 86, 194, 194, 247, 247, 250, 250, 107, 107, 253, 253, 167, 167, 181, 181, 76, 76, 261, 261, 99, 99, 266, 266, 129, 129, 269, 269, 146, 146, 89, 89, 276, 276, 102, 102, 186, 186, 98, 98, 283, 283, 163, 163, 180, 180, 60, 60, 292, 292, 42, 42, 295, 295, 297, 297, 285, 285, 109, 109, 38, 38, 305, 305, 308, 308, 119, 119, 151, 151, 49, 49, 36, 36, 309, 309, 320, 320, 182, 182, 65, 65, 196, 196, 130, 130, 179, 179, 70, 70, 190, 190, 67, 67, 80, 80, 208, 208, 164, 164, 83, 83, 345, 345, 218, 218, 128, 128, 351, 351, 353, 353, 116, 116, 358, 358, 337, 337, 85, 85, 117, 117, 366, 366, 133, 133, 168, 168, 71, 71, 373, 373, 95, 95, 211, 211, 113, 113, 249, 249, 150, 150, 385, 385, 359, 359, 177, 177, 374, 374, 394, 394, 307, 307, 398, 398, 203, 203, 401, 401, 404, 404, 406, 406, 316, 316, 409, 409, 131, 131, 414, 414, 415, 415, 78, 78, 420, 420, 275, 275, 166, 166, 426, 426, 144, 144, 430, 430, 265, 265, 254, 254, 410, 410, 438, 438, 300, 300, 105, 105, 443, 443, 357, 357, 447, 447, 29, 29, 452, 452, 453, 453, 403, 403, 458, 458, 262, 262, 206, 206, 463, 463, 171, 171, 468, 468, 284, 284, 471, 471, 159, 159, 476, 476, 306, 306, 479, 479, 482, 482, 288, 288, 56, 56, 61, 61, 79, 79, 92, 92, 101, 101, 138, 138, 140, 140, 155, 155, 162, 162, 169, 169, 170, 170, 175, 175, 184, 184, 185, 185, 189, 189, 193, 193, 195, 195, 200, 200, 209, 209, 213, 213, 214, 214, 224, 224, 226, 226, 229, 229, 233, 233, 235, 235, 240, 240, 248, 248, 270, 270, 286, 286, 287, 287, 291, 291, 293, 293, 294, 294, 296, 296, 298, 298, 299, 299, 310, 310, 315, 315, 317, 317, 318, 318, 319, 319, 321, 321, 322, 322, 325, 325, 326, 326, 329, 329, 330, 330, 333, 333, 334, 334, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 346, 346, 352, 352, 354, 354, 360, 360, 365, 365, 369, 369, 370, 370, 375, 375, 376, 376, 386, 386, 393, 393, 397, 397, 399, 399, 400, 400, 402, 402, 405, 405, 411, 411, 412, 412, 413, 413, 416, 416, 419, 419, 421, 421, 422, 422, 425, 425, 429, 429, 437, 437, 444, 444, 445, 445, 446, 446, 448, 448, 451, 451, 454, 454, 455, 455, 456, 456, 457, 457, 464, 464, 465, 465, 466, 466, 467, 467, 469, 469, 470, 470, 472, 472, 475, 475, 477, 477, 478, 478, 480, 480, 481, 481, 483, 483, 484, 484, 487, 487, 488, 488, 489, 489, 490, 490, 491, 491, 492, 492, 497, 497, 498, 498, 503, 503, 504, 504, 509, 509, 510, 510, 511, 511, 512, 512, 517, 517, 518, 518, 523, 523, 524, 524, 529, 529, 530, 530, 535, 535, 536, 536, 541, 541, 542, 542, 549, 549, 550, 550, 555, 555, 556, 556, 557, 557, 558, 558, 561, 561, 562, 562, 563, 563, 564, 564, 565, 565, 566, 566, 567, 567, 568, 568, 569, 569, 570, 570, 575, 575, 576, 576, 577, 577, 578, 578, 603, 603, 604, 604, 623, 623, 624, 624, 625, 625, 626, 626, 627, 627, 628, 628, 629, 629, 630, 630, 637, 637, 638, 638, 641, 641, 642, 642, 653, 653, 654, 654, 661, 661, 662, 662, 663, 663, 664, 664, 665, 665, 666, 666, 667, 667, 668, 668, 671, 671, 672, 672, 677, 677, 678, 678, 679, 679, 680, 680, 681, 681, 682, 682, 685, 685, 686, 686, 687, 687, 688, 688, 689, 689, 690, 690, 691, 691, 692, 692, 693, 693, 694, 694, 695, 695, 696, 696, 697, 697, 698, 698, 699, 699, 700, 700, 701, 701, 702, 702, 715, 715, 716, 716, 717, 717, 718, 718, 727, 727, 728, 728, 729, 729, 730, 730, 751, 751, 752, 752, 753, 753, 754, 754, 759, 759, 760, 760, 761, 761, 762, 762, 763, 763, 764, 764, 765, 765, 766, 766, 791, 791, 792, 792, 793, 793, 794, 794, 803, 803, 804, 804, 805, 805, 806, 806, 819, 819, 820, 820, 821, 821, 822, 822, 823, 823, 824, 824, 825, 825, 826, 826, 839, 839, 840, 840, 841, 841, 842, 842, 851, 851, 852, 852, 853, 853, 854, 854, 863, 863, 864, 864, 865, 865, 866, 866, 867, 867, 868, 868, 869, 869, 870, 870, 943, 943, 944, 944, 945, 945, 946, 946, 947, 947, 948, 948, 949, 949, 950, 950, 975, 975, 976, 976, 977, 977, 978, 978, 979, 979, 980, 980, 981, 981, 982, 982),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10, 5, 5, 6, 6, 7, 7, 8, 8, 11, 11, 12, 12, 13, 13, 14, 14, 15, 15, 16, 16, 17, 17, 18, 18, 19, 19, 20, 20, 21, 21, 22, 22, 23, 23, 24, 24, 25, 25, 26, 26, 27, 27, 28, 28, 29, 29, 30, 30, 31, 31, 32, 32, 33, 33, 34, 34, 35, 35, 36, 36, 37, 37, 38, 38, 39, 39, 40, 40, 41, 41, 42, 42, 43, 43, 44, 44, 45, 45, 46, 46, 47, 47, 48, 48, 49, 49, 50, 50, 51, 51, 52, 52, 53, 53, 54, 54, 55, 55, 56, 56, 57, 57, 58, 58, 59, 59, 60, 60, 61, 61, 62, 62, 63, 63, 64, 64, 65, 65, 66, 66, 67, 67, 68, 68, 69, 69, 70, 70, 71, 71, 72, 72, 73, 73, 74, 74, 75, 75, 76, 76, 77, 77, 78, 78, 79, 79, 80, 80, 81, 81, 82, 82, 83, 83, 84, 84, 85, 85, 86, 86, 87, 87, 88, 88, 89, 89, 90, 90, 91, 91, 92, 92, 93, 93, 94, 94, 95, 95, 96, 96, 97, 97, 98, 98, 99, 99, 100, 100, 101, 101, 102, 102, 103, 103, 104, 104, 105, 105, 106, 106, 107, 107, 108, 108, 109, 109, 110, 110, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 117, 117, 118, 118, 119, 119, 120, 120, 121, 121, 122, 122, 123, 123, 124, 124, 125, 125, 126, 126, 127, 127, 128, 128, 129, 129, 130, 130, 131, 131, 132, 132, 133, 133, 134, 134, 135, 135, 136, 136, 137, 137, 138, 138, 139, 139, 140, 140, 141, 141, 142, 142, 143, 143, 144, 144, 145, 145, 146, 146, 147, 147, 148, 148, 149, 149, 150, 150, 151, 151, 152, 152, 153, 153, 154, 154, 155, 155, 156, 156, 157, 157, 158, 158, 159, 159, 160, 160, 161, 161, 162, 162, 163, 163, 164, 164, 165, 165, 166, 166, 167, 167, 168, 168, 169, 169, 170, 170, 171, 171, 172, 172, 173, 173, 174, 174, 175, 175, 176, 176, 177, 177, 178, 178, 179, 179, 180, 180, 181, 181, 182, 182, 183, 183, 184, 184, 185, 185, 186, 186, 187, 187, 188, 188, 189, 189, 190, 190, 191, 191, 192, 192, 193, 193, 194, 194, 195, 195, 196, 196, 197, 197, 198, 198, 199, 199, 200, 200, 201, 201, 202, 202, 203, 203, 204, 204, 205, 205, 206, 206, 207, 207, 208, 208, 209, 209, 210, 210, 211, 211, 212, 212, 213, 213, 214, 214, 215, 215, 216, 216, 217, 217, 218, 218, 219, 219, 220, 220, 221, 221, 222, 222, 223, 223, 224, 224, 225, 225, 226, 226, 227, 227, 228, 228, 229, 229, 230, 230, 231, 231, 232, 232, 233, 233, 234, 234, 235, 235, 236, 236, 237, 237, 238, 238, 239, 239, 240, 240, 241, 241, 242, 242, 243, 243, 244, 244, 245, 245, 246, 246, 247, 247, 248, 248, 249, 249, 250, 250, 251, 251, 252, 252, 253, 253, 254, 254, 255, 255, 256, 256, 257, 257, 258, 258, 259, 259, 260, 260, 261, 261, 262, 262, 263, 263, 264, 264, 265, 265, 266, 266, 267, 267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 272, 273, 273, 274, 274, 275, 275, 276, 276, 277, 277, 278, 278, 279, 279, 280, 280, 281, 281, 282, 282, 283, 283, 284, 284, 285, 285, 286, 286, 287, 287, 288, 288, 289, 289, 290, 290, 291, 291, 292, 292, 293, 293, 294, 294, 295, 295, 296, 296, 297, 297, 298, 298, 299, 299, 300, 300, 301, 301, 302, 302, 303, 303, 304, 304, 305, 305, 306, 306, 307, 307, 308, 308, 309, 309, 310, 310, 311, 311, 312, 312, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 323, 323, 324, 324, 325, 325, 326, 326, 327, 327, 328, 328, 329, 329, 330, 330, 331, 331, 332, 332, 333, 333, 334, 334, 335, 335, 336, 336, 337, 337, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 345, 345, 346, 346, 347, 347, 348, 348, 349, 349, 350, 350, 351, 351, 352, 352, 353, 353, 354, 354, 355, 355, 356, 356, 357, 357, 358, 358, 359, 359, 360, 360, 361, 361, 362, 362, 363, 363, 364, 364, 365, 365, 366, 366, 367, 367, 368, 368, 369, 369, 370, 370, 371, 371, 372, 372, 373, 373, 374, 374, 375, 375, 376, 376, 377, 377, 378, 378, 379, 379, 380, 380, 381, 381, 382, 382, 383, 383, 384, 384, 385, 385, 386, 386, 387, 387, 388, 388, 389, 389, 390, 390, 391, 391, 392, 392, 393, 393, 394, 394, 395, 395, 396, 396, 397, 397, 398, 398, 399, 399, 400, 400, 401, 401, 402, 402, 403, 403, 404, 404, 405, 405, 406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 412, 412, 413, 413, 414, 414, 415, 415, 416, 416, 417, 417, 418, 418, 419, 419, 420, 420, 421, 421, 422, 422, 423, 423, 424, 424, 425, 425, 426, 426, 427, 427, 428, 428, 429, 429, 430, 430, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446, 447, 447, 448, 448, 449, 449, 450, 450, 451, 451, 452, 452, 453, 453, 454, 454, 455, 455, 456, 456, 457, 457, 458, 458, 459, 459, 460, 460, 461, 461, 462, 462, 463, 463, 464, 464, 465, 465, 466, 466, 467, 467, 468, 468, 469, 469, 470, 470, 471, 471, 472, 472, 473, 473, 474, 474, 475, 475, 476, 476, 477, 477, 478, 478, 479, 479, 480, 480, 481, 481, 482, 482, 483, 483, 484, 484, 485, 485, 486, 486, 487, 487, 488, 488, 489, 489, 490, 490, 491, 491, 492, 492, 493, 493, 494, 494, 495, 495, 496, 496, 497, 497, 498, 498, 499, 499, 500, 500, 501, 501, 502, 502, 503, 503, 504, 504, 505, 505, 506, 506, 507, 507, 508, 508, 509, 509, 510, 510)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 5, 5, 3, 3, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 4, 4, 5, 5, 6, 6, 3, 3, 4, 4, 5, 5, 6, 6, 6, 6, 7, 7, 6, 6, 5, 5, 6, 6, 6, 6, 5, 5, 6, 6, 7, 7, 7, 7, 5, 5, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 4, 4, 5, 5, 6, 6, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 9, 9, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 6, 6, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 3, 3, 4, 4, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 4, 4, 5, 5, 5, 5, 6, 6, 3, 3, 4, 4, 5, 5, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 5, 5, 6, 6, 6, 6, 6, 6, 7, 7, 5, 5, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 7, 7, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 6, 6, 7, 7, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 6, 6, 8, 8, 9, 9, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 4, 4, 5, 5, 6, 6, 9, 9, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 9, 9, 7, 7, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 5, 5, 6, 6, 7, 7, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((135, 136, 141, 142, 149, 150, 155, 156, 157, 158, 161, 162, 167, 168, 173, 174, 175, 176, 187, 188, 189, 190, 195, 196, 203, 204, 205, 206, 211, 212, 219, 220, 223, 224, 225, 226, 231, 232, 235, 236, 257, 258, 267, 268, 275, 276, 281, 282, 287, 288, 293, 294, 301, 302, 305, 306, 315, 316, 319, 320, 321, 322, 323, 324, 337, 338, 339, 340, 341, 342, 349, 350, 351, 352, 359, 360, 361, 362, 363, 364, 371, 372, 383, 384, 385, 386, 389, 390, 391, 392, 405, 406, 409, 410, 425, 426, 447, 448, 449, 450, 459, 460, 463, 464, 467, 468, 473, 474, 475, 476, 477, 478, 479, 480, 485, 486, 487, 488, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 505, 506, 507, 508, 513, 514, 517, 518, 519, 520, 523, 524, 525, 526, 527, 528, 531, 532, 533, 534, 535, 536, 541, 542, 543, 544, 547, 548, 551, 552, 555, 556, 557, 558, 559, 560, 565, 566, 567, 568, 569, 570, 575, 576, 577, 578, 579, 580, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 609, 610, 611, 612, 617, 618, 619, 620, 625, 626, 631, 632, 633, 634, 635, 636, 637, 638, 643, 644, 645, 646, 649, 650, 651, 652, 653, 654, 657, 658, 659, 660, 669, 670, 671, 672, 673, 674, 677, 678, 679, 680, 683, 684, 685, 686, 689, 690, 691, 692, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725, 726, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 839, 840, 841, 842, 847, 848, 849, 850, 855, 856, 857, 858, 863, 864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (121, 122, 125, 126, 135, 136, 141, 142, 147, 148, 153, 154, 157, 158, 187, 188, 191, 192, 197, 198, 201, 202, 215, 216, 219, 220, 221, 222, 227, 228, 231, 232, 237, 238, 241, 242, 243, 244, 245, 246, 251, 252, 255, 256, 257, 258, 259, 260, 263, 264, 267, 268, 271, 272, 273, 274, 277, 278, 279, 280, 281, 282, 289, 290, 301, 302, 303, 304, 311, 312, 313, 314, 323, 324, 327, 328, 331, 332, 335, 336, 347, 348, 349, 350, 355, 356, 361, 362, 363, 364, 367, 368, 371, 372, 377, 378, 379, 380, 381, 382, 383, 384, 387, 388, 389, 390, 391, 392, 395, 396, 407, 408, 417, 418, 423, 424, 427, 428, 431, 432, 433, 434, 435, 436, 439, 440, 441, 442, 449, 450, 459, 460, 461, 462, 473, 474, 485, 486, 493, 494, 495, 496, 499, 500, 501, 502, 505, 506, 507, 508, 513, 514, 515, 516, 519, 520, 521, 522, 525, 526, 527, 528, 531, 532, 533, 534, 537, 538, 539, 540, 543, 544, 545, 546, 547, 548, 551, 552, 553, 554, 559, 560, 571, 572, 573, 574, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 631, 632, 633, 634, 635, 636, 639, 640, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 655, 656, 657, 658, 659, 660, 669, 670, 673, 674, 675, 676, 683, 684, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 719, 720, 721, 722, 723, 724, 725, 726, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 755, 756, 757, 758, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 795, 796, 797, 798, 799, 800, 801, 802, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 843, 844, 845, 846, 847, 848, 849, 850, 855, 856, 857, 858, 859, 860, 861, 862, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 759, 760, 761, 762, 763, 764, 765, 766, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 863, 864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 1, 1, 1, 2, 1, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 2, 0, 1, 1, 1, 2, 0, 0, 1, 0, 1, 2, 1, 2, 0, 0, 0, 2, 2, -2, 0, 0, 1, 1, 2, 1, 1, 1, 1, 2, 0, -2, -2, -2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 1, 2, 0, 0, 0, 2, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 1, -2, 0, 0, 1, 1, 0, 1, 2, -2, 0, -2, 1, 1, 0, -2, 2, 2, 0, 2, -2, -2, 1, 2, 0, 2, 0, 0, -2, -2, 0, -2, -2, 2, -2, 1, 0, -2, 1, -2, 1, 1, 1, 2, 0, 0, 0, 1, 2, -2, -2, 1, -2, -2, 0, 0, 0, 2, 2, 0, -2, -2, 0, 0, 1, -2, 0, 0, 0, 1, -2, -2, 1, 0, 1, 1, 0, -2, 1, 0, -2, 0, -2, -2, 2, -2, -2, -2, 0, -2, -2, -2, 0, -2, 1, 1, -2, -2, 1, 0, -2, 2, 0, 2, -2, -2, -2, 1, -2, 0, -2, -2, -2, 2, -2, -2, -2, -2, -2, 2, -2, -2, 1, 2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, -2, 1, -2, -2, -2, 1, -2, -2, -2, -2, 2, -2, 1, -2, -2, -2, -2, -2, -2, 0, 0, 0, 2, -2, 2, -2, -2, -2, -2, -2, -2, 2, 0, 1, 1, -2, -2, -2, -2, 1, 1, 1, 2, 0, 2, -2, 1, -2, -2, 1, -2, -2, -2, -2, 2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, -2, 1, -2, -2, -2, -2, -2, 1, -2, -2, -2, -2, 0, -2, 1, -2, -2, -2, -2, 2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, 2, 0, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, 0, -2, -2, -2, 2, 1, -2, 1, -2, -2, -2, -2, -2, -2, 0, 2, -2, 0, -2, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, -2, 0, 1, -2, -2, 2, -2, -2, -2, -2, 0, -2, -2, -2, 0, -2, -2, 1, -2, -2, 2, -2, -2, -2, 0, -2, -2, 0, -2, -2, -2, -2, 0, -2, 1, 1, -2, -2, -2, -2, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 2, 2, 1, 1, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, 1, 0, 2, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, 0, 1, 2, 0, 2, 2, 2, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, -2, 1, 1, 1, 0, 0, -2, 1, 1, -2, 0, 2, -2, 0, 0, 0, 2, 0, 1, 1, 1, 2, 1, 0, -2, -2, 2, 1, 0, 0, 1, 1, 2, 1, -2, 0, 1, 2, 0, 1, 0, -2, 2, 0, 0, 0, 1, 0, -2, -2, 0, -2, -2, -2, -2, -2, 1, 2, 0, -2, 0, -2, -2, -2, 1, 2, -2, 0, -2, -2, -2, -2, 0, 1, 1, 1, -2, -2, 2, -2, 1, 2, 0, -2, -2, -2, 1, 2, 1, 0, 0, 0, 1, 1, 0, 1, -2, -2, -2, 1, 1, -2, -2, -2, 0, -2, 1, 1, -2, -2, 0, 2, 0, 0, 0, -2, 1, 1, 2, 2, 1, 0, -2, 2, -2, -2, 1, -2, -2, 1, 2, -2, -2, -2, -2, 1, 0, 2, -2, 2, -2, 1, -2, -2, 2, 2, 0, 0, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, 1, 0, 1, 2, 1, -2, -2, -2, 2, 0, -2, -2, 1, 1, -2, -2, -2, -2, 1, 0, 1, -2, -2, -2, 0, 0, 2, 0, 0, 0, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, 2, -2, 1, -2, -2, 1, 2, -2, -2, -2, 1, -2, -2, -2, -2, -2, 1, -2, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, 1, -2, -2, 2, -2, -2, -2, 2, -2, -2, -2, 0, 0, 1, 2, -2, -2, 0, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, 1, -2, -2, 0, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, 1, 0, -2, -2, -2, 2, 0, -2, -2, -2, 1, -2, -2, -2, -2, 1, -2, 1, -2, -2, 0, -2, 0, 2, 1, 1, -2, -2, -2, -2, 0, -2, -2, -2, -2, -2, 1, 1, -2, -2, -2, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2, 0, -2, -2, 1, -2, -2, -2, -2, 2, -2, -2, 1, 0, -2, 2, 1, -2, -2, -2, -2, 0, -2, -2, -2, 1, -2, -2, -2, -2, -2, 1, -2, 2, 0, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, 1, -2, -2, -2, 1, -2, -2, 0, -2, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 0, 0, -2, -2, -2, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((143257, 6999, 220619, 35159, 102496, 2865, 4936, 11682, 296115, 10141, 536, 9457, 3798, 8137, 9405, 438, 11162, 874, 10905, 12264, 188370, 9170, 438, 189082, 168644, 41132, 60757, 536, 77449, 12703, 13359, 7856, 536, 112477, 128407, 12213, 343001, 11768, 438, 13341, 536, 163298, 169876, 178654, 366, 536, -1024, 138400, 113147, 10063, 10426, 536, 11583, 10911, 11135, 13214, 655, 2509, -1024, -1024, -1024, 56288, 6053, 6073, 87936, 210259, 14325, 21588, 31288, 17574, 536, 10599, 11358, 254835, 282656, 12740, 366, 280953, 274352, 61379, 536, 72176, 63306, 72768, 8933, 62681, 536, 100812, 7841, 1913, 2634, 1379, -1024, 43861, 55801, 5452, 5884, 122124, 8833, 366, -1024, 256505, -1024, 13924, 14280, 243041, -1024, 655, 655, 120570, 655, -1024, -1024, 8696, 366, 174854, 438, 173562, 191652, -1024, -1024, 201552, -1024, -1024, 655, -1024, 13187, 30576, -1024, 3304, -1024, 7101, 7450, 10849, 366, 258917, 229344, 238128, 11957, 366, -1024, -1024, 7426, -1024, -1024, 199641, 219728, 194686, 438, 366, 207613, -1024, -1024, 122647, 106823, 8440, -1024, 105754, 115313, 86370, 7181, -1024, -1024, 13918, 215126, 11857, 12086, 155417, -1024, 2257, 17765, -1024, 23247, -1024, -1024, 655, -1024, -1024, -1024, 198683, -1024, -1024, -1024, 168345, -1024, 9550, 10000, -1024, -1024, 4009, 46551, -1024, 438, 40205, 536, -1024, -1024, -1024, 5356, -1024, 56600, -1024, -1024, -1024, 655, -1024, -1024, -1024, -1024, -1024, 366, -1024, -1024, 13457, 366, -1024, 14134, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 655, -1024, -1024, 12661, -1024, -1024, -1024, 12117, -1024, -1024, -1024, -1024, 366, -1024, 10717, -1024, -1024, -1024, -1024, -1024, -1024, 86721, 93271, 79360, 536, -1024, 655, -1024, -1024, -1024, -1024, -1024, -1024, 366, 92619, 6353, 6881, -1024, -1024, -1024, -1024, 13519, 14365, 13074, 366, 327188, 438, -1024, 14116, -1024, -1024, 8458, -1024, -1024, -1024, -1024, 438, -1024, -1024, -1024, 266292, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 179309, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 655, -1024, 7422, -1024, -1024, -1024, -1024, -1024, 8558, -1024, -1024, -1024, -1024, 309503, -1024, 14051, -1024, -1024, -1024, -1024, 438, -1024, 142036, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 366, 240415, -1024, 11414, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 17594, -1024, -1024, -1024, 4462, -1024, -1024, -1024, 202264, -1024, -1024, -1024, 366, 13231, -1024, 13141, -1024, -1024, -1024, -1024, -1024, -1024, 159694, 366, -1024, 150454, -1024, -1024, -1024, -1024, -1024, 13422, -1024, -1024, -1024, 8717, -1024, -1024, -1024, 174286, 11616, -1024, -1024, 536, -1024, -1024, -1024, -1024, 219896, -1024, -1024, -1024, 19133, -1024, -1024, 4482, -1024, -1024, 536, -1024, -1024, -1024, 81014, -1024, -1024, 92288, -1024, -1024, -1024, -1024, 93549, -1024, 9373, 9224, -1024, -1024, -1024, -1024, 360863, 366, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024),
                (174607, 6556, 255008, 45076, 123069, 2859, 67804, 11180, 311672, 10141, 536, 8405, 9521, 366, 536, 12369, 13164, 12800, 25512, 1027, 2278, 5161, 6200, 4772, 536, 9964, 11486, 136920, 167478, 12829, 210031, 655, 221268, 12716, 342909, 12093, 438, 13085, 267279, 87202, 106721, 62499, 438, 6915, 536, 8246, 8861, 128609, 147650, 9350, 366, 212188, 438, 438, 438, 231170, 194134, 184262, 207596, 10236, 236101, 655, 11032, 62222, 55491, 24565, 4013, 33263, 4621, 2665, 9979, -1024, 879, 13465, 14728, 101641, 109524, -1024, 8957, 5556, -1024, 219629, 366, -1024, 50623, 14659, 19800, 536, 22897, 3458, 3954, 2944, 536, 11560, 245448, -1024, -1024, 438, 10438, 164029, 133235, 12000, 13030, 655, 13357, -1024, 156749, 6635, 536, 86298, 7796, 70949, -1024, 366, 292223, 299755, 269333, 9968, 128963, -1024, -1024, 189047, -1024, -1024, -1024, -1024, -1024, 11613, 366, 291503, -1024, 278829, -1024, -1024, -1024, 7255, 366, -1024, 150501, -1024, -1024, -1024, -1024, 97284, 8182, 7315, 8138, -1024, -1024, 655, -1024, 4206, 438, 58980, -1024, -1024, -1024, 5367, 438, 5517, 65864, 250490, 245723, 12901, 13128, 212371, 13212, -1024, -1024, -1024, 13938, 14002, -1024, -1024, -1024, 202296, -1024, 10798, 11122, -1024, -1024, 128086, 438, 145844, 127495, 137881, -1024, 9219, 9605, 536, 655, 8857, 108228, -1024, 366, -1024, -1024, 10664, -1024, -1024, 10910, 366, -1024, -1024, -1024, -1024, 1632, 10512, 655, -1024, 366, -1024, 13968, -1024, -1024, 536, 655, 40898, 33271, -1024, -1024, -1024, -1024, -1024, 147674, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 7676, -1024, -1024, 13243, 353140, 12782, 366, 13655, -1024, -1024, -1024, 655, 159960, -1024, -1024, 10526, 10864, -1024, -1024, -1024, -1024, 12691, 196896, 13023, -1024, -1024, -1024, 71564, 82374, 366, 89600, 79702, 72123, -1024, -1024, -1024, -1024, -1024, -1024, 7692, -1024, -1024, -1024, 536, -1024, 13437, -1024, -1024, 14343, 366, -1024, -1024, -1024, 11898, -1024, -1024, -1024, -1024, -1024, 13380, -1024, 366, 11785, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 284139, -1024, 8238, -1024, -1024, 655, -1024, -1024, -1024, 438, -1024, -1024, -1024, 169081, 174546, 10051, 366, -1024, -1024, 194459, -1024, -1024, -1024, 178275, -1024, -1024, -1024, -1024, -1024, -1024, 327333, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 5605, 5964, -1024, -1024, 55753, -1024, -1024, -1024, -1024, 38714, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 10791, 174578, -1024, -1024, -1024, 366, 54302, -1024, -1024, -1024, 8400, -1024, -1024, -1024, -1024, 10398, -1024, 10857, -1024, -1024, 92392, -1024, 81259, 655, 8536, 8924, -1024, -1024, -1024, -1024, 87409, -1024, -1024, -1024, -1024, -1024, 2930, 3492, -1024, -1024, -1024, 366, 324470, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, 86584, -1024, -1024, 2916, -1024, -1024, -1024, -1024, 655, -1024, -1024, 13684, 360960, -1024, 366, 14100, -1024, -1024, -1024, -1024, 250736, -1024, -1024, -1024, 12731, -1024, -1024, -1024, -1024, -1024, 9356, -1024, 366, 194726, -1024, -1024, -1024, 55835, -1024, -1024, -1024, -1024, -1024, -1024, 5985, -1024, -1024, -1024, 11628, -1024, -1024, 360032, -1024, -1024, 497, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024),
                (270729, 6667, 360960, 67917, 148442, -1024, -1024, -1024, -1024, 12327, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024, -1024)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((154, 73, 167, 132, 17, 56, 158, 137, 170, 162, 38, 119, 10, 4, 51, 129, 14, 27, 155, 6, 86, 169, 111, 46, 152, 169, 130, 31, 159, 50, 140, 84, 160, 153, 35, 160, 170, 169, 109, 36, 159, 110, 19, 9, 98, 39, 0, 3, 94, 25, 124, 106, 168, 31, 152, 168, 92, 85, 0, 0, 171, 7, 71, 127, 168, 43, 161, 43, 1, 3, 128, 46, 142, 59, 9, 18, 91, 39, 143, 159, 92, 37, 156, 21, 1, 2, 73, 29, 156, 107, 165, 158, 0, 110, 21, 39, 161, 7, 89, 146, 0, 132, 171, 83, 164, 118, 0, 66, 148, 160, 82, 32, 144, 170, 151, 94, 162, 11, 155, 0, 171, 109, 0, 0, 49, 0, 102, 85, 171, 34, 171, 18, 107, 170, 147, 78, 169, 14, 142, 93, 171, 0, 146, 171, 66, 28, 1, 6, 94, 19, 155, 9, 85, 134, 169, 100, 171, 158, 31, 85, 7, 0, 171, 19, 114, 26, 105, 85, 0, 169, 120, 0, 158, 0, 137, 76, 0, 0, 137, 157, 68, 171, 43, 142, 171, 85, 166, 10, 78, 153, 170, 171, 66, 16, 146, 114, 0, 0, 46, 171, 14, 91, 155, 171, 114, 57, 171, 85, 0, 85, 164, 85, 0, 2, 40, 0, 85, 171, 34, 85, 171, 171, 57, 137, 62, 171, 102, 171, 119, 43, 171, 39, 0, 27, 114, 122, 171, 171, 57, 0, 34, 0, 68, 114, 0, 123, 171, 171, 85, 9, 0, 1, 57, 0, 146, 102, 171, 0, 68, 128, 171, 156, 170, 105, 168, 171, 28, 122, 171, 168, 171, 170, 138, 19, 166, 0, 51, 102, 0, 114, 171, 171, 57, 0, 34, 0, 85, 171, 137, 57, 171, 133, 171, 171, 114, 171, 114, 171, 114, 43, 0, 171, 114, 0, 57, 133, 171, 114, 171, 0, 57, 57, 0, 114, 171, 0, 57, 0, 15, 0, 85, 0, 57, 171, 114, 0, 26, 68, 0, 114, 163, 154, 171, 98, 171, 57, 128, 0, 19, 0, 49, 85, 0, 171, 114, 114, 171, 137, 171, 171, 165, 146, 171, 78, 171, 107, 0, 128, 171, 114, 57, 171, 156, 102, 171, 0, 13, 85, 0, 171, 146, 114, 171, 171, 164, 114, 171, 142, 57, 114, 171, 85, 122, 171, 166, 146, 171, 85, 171, 57, 102, 28, 4, 19, 0, 0, 57, 156, 171, 171, 114, 169, 155, 114, 171, 158, 171, 114, 171, 0, 11, 57, 0, 0, 13, 57, 0, 167, 171, 171, 114, 57, 171, 0, 8, 57, 0, 164, 171, 171, 114, 0, 2, 57, 1, 19, 0, 0, 57, 171, 170, 114, 171, 0, 171, 0, 0, 0, 0, 0, 0, 171, 171, 0, 0, 0, 0, 171, 171, 0, 0, 0, 0, 171, 171, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 0, 0, 171, 171, 0, 0, 0, 0, 0, 0, 68, 68, 171, 171, 43, 43, 171, 171, 171, 171, 0, 0, 171, 171, 171, 171, 85, 85, 0, 0, 85, 85, 171, 171, 171, 171, 102, 102, 171, 171, 43, 43, 171, 171, 0, 0, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 102, 102, 0, 0, 171, 171, 0, 0, 0, 0, 85, 85, 171, 171, 171, 171, 114, 114, 0, 0, 57, 57, 171, 171, 0, 0, 57, 57, 114, 114, 171, 171, 0, 0, 57, 57, 0, 0, 0, 0, 0, 0, 57, 57, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 114, 114, 171, 171, 137, 137, 171, 171, 171, 171, 171, 171, 171, 171, 114, 114, 57, 57, 171, 171, 0, 0, 85, 85, 0, 0, 171, 171, 114, 114, 171, 171, 171, 171, 171, 171, 57, 57, 171, 171, 171, 171, 171, 171, 0, 0, 171, 171, 171, 171, 114, 114, 114, 114, 171, 171, 171, 171, 0, 0, 57, 57, 0, 0, 0, 0, 57, 57, 0, 0, 171, 171, 171, 171, 57, 57, 171, 171, 0, 0, 57, 57, 0, 0, 171, 171, 0, 0, 57, 57, 0, 0, 171, 171, 171, 171, 0, 0, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 137, 137, 137, 137, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 85, 85, 85, 85, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 57, 57, 57, 57, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 57, 57, 57, 57, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171),
                (137, 50, 165, 115, 17, 38, 161, 130, 169, 167, 50, 6, 53, 149, 21, 19, 128, 93, 11, 25, 158, 126, 169, 166, 37, 5, 50, 134, 14, 164, 90, 39, 154, 157, 170, 169, 88, 19, 165, 22, 2, 5, 92, 39, 147, 100, 164, 160, 47, 170, 134, 47, 161, 48, 7, 24, 116, 24, 159, 4, 130, 78, 159, 15, 98, 1, 31, 124, 8, 69, 8, 0, 153, 6, 99, 128, 24, 0, 101, 50, 171, 9, 75, 171, 9, 170, 121, 21, 159, 88, 165, 159, 34, 46, 155, 124, 0, 39, 2, 10, 114, 7, 52, 111, 6, 171, 53, 0, 23, 1, 71, 123, 0, 66, 9, 18, 142, 44, 126, 171, 16, 123, 0, 62, 171, 68, 156, 171, 143, 70, 171, 19, 171, 10, 171, 9, 68, 0, 141, 51, 158, 32, 133, 117, 164, 43, 147, 171, 0, 108, 171, 169, 121, 71, 171, 0, 171, 4, 55, 27, 142, 0, 20, 13, 102, 49, 1, 0, 94, 171, 43, 71, 171, 122, 0, 138, 171, 85, 166, 76, 171, 169, 143, 89, 167, 14, 171, 0, 9, 47, 1, 9, 158, 0, 85, 0, 171, 85, 171, 171, 28, 73, 171, 0, 171, 0, 39, 146, 7, 0, 33, 0, 96, 149, 43, 33, 2, 14, 102, 0, 171, 0, 95, 171, 131, 78, 162, 57, 171, 163, 85, 171, 98, 0, 171, 166, 171, 170, 118, 14, 171, 114, 11, 29, 3, 0, 70, 57, 128, 128, 21, 0, 85, 169, 137, 76, 171, 0, 137, 170, 156, 85, 169, 21, 137, 57, 171, 0, 57, 0, 85, 119, 171, 171, 0, 145, 171, 102, 171, 171, 78, 119, 171, 0, 171, 124, 171, 171, 43, 107, 171, 47, 0, 4, 30, 61, 0, 85, 0, 171, 85, 39, 3, 0, 57, 171, 139, 68, 171, 122, 171, 85, 171, 26, 0, 0, 76, 13, 0, 3, 95, 0, 171, 38, 0, 0, 114, 43, 0, 0, 73, 171, 114, 0, 64, 102, 0, 171, 114, 1, 20, 114, 171, 98, 43, 0, 57, 128, 171, 171, 114, 128, 171, 43, 0, 0, 43, 0, 57, 158, 171, 171, 68, 21, 0, 0, 114, 0, 13, 0, 73, 171, 114, 171, 114, 57, 0, 34, 0, 0, 28, 57, 0, 171, 161, 114, 171, 68, 171, 158, 171, 171, 102, 0, 7, 102, 2, 28, 0, 3, 0, 1, 23, 4, 146, 43, 0, 171, 114, 149, 171, 171, 114, 0, 28, 0, 10, 85, 0, 171, 162, 137, 171, 57, 171, 19, 0, 0, 9, 0, 14, 57, 0, 12, 0, 0, 57, 0, 6, 0, 38, 169, 171, 171, 132, 64, 171, 102, 0, 0, 9, 57, 0, 171, 161, 114, 171, 9, 0, 171, 168, 114, 169, 160, 171, 102, 171, 5, 0, 0, 57, 3, 0, 171, 168, 114, 171, 171, 168, 114, 171, 170, 171, 171, 142, 114, 171, 57, 57, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 171, 171, 171, 171, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 171, 171, 57, 57, 171, 171, 171, 171, 171, 171, 0, 0, 85, 85, 171, 171, 0, 0, 137, 137, 57, 57, 171, 171, 0, 0, 85, 85, 171, 171, 171, 171, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 171, 171, 114, 114, 0, 0, 171, 171, 114, 114, 128, 128, 171, 171, 128, 128, 171, 171, 43, 43, 0, 0, 0, 0, 57, 57, 171, 171, 68, 68, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 102, 102, 0, 0, 102, 102, 0, 0, 171, 171, 171, 171, 114, 114, 85, 85, 0, 0, 171, 171, 171, 171, 57, 57, 171, 171, 0, 0, 0, 0, 0, 0, 57, 57, 0, 0, 171, 171, 171, 171, 102, 102, 0, 0, 0, 0, 57, 57, 0, 0, 171, 171, 114, 114, 171, 171, 171, 171, 114, 114, 171, 171, 102, 102, 171, 171, 0, 0, 0, 0, 57, 57, 171, 171, 114, 114, 171, 171, 171, 171, 114, 114, 171, 171, 171, 171, 171, 171, 114, 114, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 128, 128, 128, 128, 171, 171, 171, 171, 43, 43, 43, 43, 0, 0, 0, 0, 171, 171, 171, 171, 68, 68, 68, 68, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 85, 85, 85, 85, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 114, 114, 114, 114, 171, 171, 171, 171, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 114, 114, 114, 114, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 0, 0, 0, 0, 0, 0, 0, 0, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 114, 114, 114, 114, 114, 114, 114, 114, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171),
                (85, 27, 167, 79, 12, 22, 166, 3, 39, 145, 171, 170, 76, 22, 22, 166, 166, 3, 3, 39, 39, 171, 171, 170, 170, 76, 76, 22, 22, 22, 22, 166, 166, 166, 166, 3, 3, 3, 3, 39, 39, 39, 39, 171, 171, 171, 171, 170, 170, 170, 170, 76, 76, 76, 76, 22, 22, 22, 22, 22, 22, 22, 22, 166, 166, 166, 166, 166, 166, 166, 166, 3, 3, 3, 3, 3, 3, 3, 3, 39, 39, 39, 39, 39, 39, 39, 39, 171, 171, 171, 171, 171, 171, 171, 171, 170, 170, 170, 170, 170, 170, 170, 170, 76, 76, 76, 76, 76, 76, 76, 76, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 7, 5, 13, 11, 25, 9, 35, 21, 19, 17, 67, 83, 15, 31, 45, 57, 89, 145, 29, 113, 23, 43, 51, 189, 27, 61, 63, 41, 55, 33, 153, 139, 97, 37, 269, 133, 39, 73, 101, 107, 123, 239, 71, 47, 445, 337, 49, 175, 109, 53, 401, 167, 203, 369, 65, 59, 447, 449, 451, 197, 93, 79, 261, 163, 301, 69, 365, 413, 127, 121, 179, 75, 213, 231, 77, 151, 245, 209, 81, 187, 329, 85, 249, 317, 87, 131, 227, 91, 169, 225, 453, 95, 119, 207, 297, 325, 99, 255, 455, 103, 457, 105, 287, 201, 459, 165, 235, 291, 111, -1, -1, 383, 115, 117, 183, 303, 305, 461, 463, 381, 465, 467, 125, 469, 143, 129, 471, 195, 473, 159, 181, 349, 135, 137, 347, 309, 219, 141, 475, 477, 343, -1, -1, 147, 409, 283, 149, 321, 313, -1, -1, 155, 397, 157, 479, 307, 257, 161, 391, -1, -1, 299, 221, 211, 247, 173, 481, 361, 171, 483, 357, -1, -1, 177, 485, -1, -1, 267, 487, 489, 491, 185, 493, 223, 295, -1, -1, 191, 417, 495, 193, 315, 345, -1, -1, 497, 199, 499, 311, -1, -1, 501, 205, -1, -1, -1, -1, 503, 259, -1, -1, 393, 215, 505, 217, -1, -1, 507, 509, -1, -1, -1, -1, 511, 513, 515, 229, 517, 519, 233, 521, -1, -1, 237, 523, -1, -1, 525, 241, 527, 243, -1, -1, -1, -1, -1, -1, 251, 431, 423, 253, 529, 279, -1, -1, -1, -1, -1, -1, 263, 427, 265, 293, -1, -1, -1, -1, 271, 439, 373, 273, 275, 331, 531, 277, 533, 535, 281, 537, -1, -1, 539, 285, 541, 543, 545, 289, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 547, 549, 551, 553, 323, 555, -1, -1, 557, 559, -1, -1, 561, 563, 565, 567, 569, 319, 571, 359, 573, 575, -1, -1, 577, 327, -1, -1, -1, -1, 333, 579, 335, 581, -1, -1, 583, 339, 585, 341, -1, -1, -1, -1, 587, 589, 591, 593, 595, 351, 353, 597, 355, 599, -1, -1, -1, -1, 601, 603, 605, 363, -1, -1, 607, 367, 609, 611, 613, 371, 615, 617, 619, 375, 377, 621, 379, 623, -1, -1, -1, -1, 625, 385, 387, 627, 389, 629, -1, -1, -1, -1, 395, 631, -1, -1, 399, 633, 635, 637, 405, 403, 639, 641, 407, 643, -1, -1, 645, 411, 647, 649, 651, 415, 653, 655, 419, 657, 659, 421, 661, 663, 665, 425, 667, 669, 429, 671, -1, -1, 673, 433, 675, 435, 437, 677, -1, -1, 679, 441, 443, 681, 683, 685, 687, 689, 691, 693, 695, 697, 699, 701, 703, 705, -1, -1, 707, 709, -1, -1, -1, -1, -1, -1, -1, -1, 711, 713, -1, -1, 715, 717, -1, -1, 719, 721, -1, -1, 723, 725, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 727, 729, 731, 733, 735, 737, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 739, 741, -1, -1, -1, -1, -1, -1, -1, -1, 743, 745, -1, -1, 747, 749, 751, 753, -1, -1, -1, -1, -1, -1, 755, 757, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 759, 761, 763, 765, -1, -1, -1, -1, -1, -1, 767, 769, -1, -1, 771, 773, -1, -1, -1, -1, -1, -1, 775, 777, 779, 781, 783, 785, 787, 789, -1, -1, -1, -1, -1, -1, -1, -1, 791, 793, 795, 797, 799, 801, 803, 805, -1, -1, -1, -1, 807, 809, 811, 813, -1, -1, 815, 817, 819, 821, -1, -1, -1, -1, 823, 825, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 827, 829, 831, 833, 835, 837, 839, 841, -1, -1, -1, -1, 843, 845, 847, 849, -1, -1, -1, -1, 851, 853, -1, -1, -1, -1, -1, -1, 855, 857, 859, 861, -1, -1, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, 887, 889, 891, 893, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 895, 897, 899, 901, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 903, 905, 907, 909, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, -1, -1, -1, -1, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, -1, -1, -1, -1, 951, 953, 955, 957, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 959, 961, 963, 965, -1, -1, -1, -1, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 7, 5, 11, 17, 21, 9, 33, 49, 15, 39, 13, 45, 25, 53, 29, 19, 65, 69, 85, 23, 259, 151, 63, 97, 27, 61, 101, 253, 31, 73, 149, 35, 235, 127, 37, 113, 275, 41, 187, 107, 43, 75, 143, 47, 181, 271, 77, 459, 51, 59, 175, 55, 161, 81, 57, 327, 285, 353, 197, 117, 223, 157, 79, 415, 67, 89, 215, 71, 205, 489, 231, 323, 121, 201, 135, 491, 105, 83, 493, 293, 93, 495, 413, 347, 87, 269, 281, 91, 337, 341, 133, 95, 349, -1, -1, 99, 317, 193, 137, 243, 103, 139, 377, 497, 221, 467, 109, 429, 111, 125, 499, 115, 209, 251, 227, 119, 179, -1, -1, 123, 501, -1, -1, -1, -1, 477, 129, 131, 503, 303, 505, -1, -1, 301, 141, 507, 289, -1, -1, -1, -1, 145, 305, 147, 229, -1, -1, 171, 509, 383, 153, 155, 511, 513, 515, 363, 159, 241, 373, 449, 163, 165, 169, 167, 457, -1, -1, 517, 297, 173, 519, -1, -1, 177, 521, 247, 331, -1, -1, 389, 183, 185, 351, 345, 523, 399, 189, 191, 393, 313, 309, 525, 195, -1, -1, 199, 527, 529, 375, 203, 531, -1, -1, 533, 207, 371, 355, 535, 211, 537, 213, -1, -1, 217, 367, 267, 219, -1, -1, -1, -1, 539, 225, -1, -1, 541, 543, -1, -1, 545, 233, -1, -1, 237, 441, 419, 239, 291, 547, -1, -1, 245, 339, -1, -1, 249, 299, -1, -1, 549, 551, 453, 255, 257, 553, 555, 557, 359, 261, 263, 409, 357, 265, 559, 561, -1, -1, 563, 565, 273, 567, 569, 571, 277, 573, 279, 575, 577, 343, 283, 579, -1, -1, 287, 581, -1, -1, -1, -1, 333, 583, 427, 295, -1, -1, -1, -1, -1, -1, -1, -1, 585, 487, 587, 307, -1, -1, 311, 589, -1, -1, 315, 591, -1, -1, 319, 379, 425, 321, -1, -1, 325, 593, -1, -1, 329, 595, -1, -1, 597, 599, 601, 335, -1, -1, 603, 605, -1, -1, -1, -1, -1, -1, -1, -1, 607, 609, -1, -1, 611, 613, 615, 617, -1, -1, 619, 621, 361, 473, 623, 625, 365, 627, -1, -1, 629, 369, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 471, 381, -1, -1, 631, 385, 387, 633, -1, -1, 391, 635, 637, 639, 641, 395, 643, 397, -1, -1, 401, 645, 437, 403, 405, 407, -1, -1, -1, -1, 411, 647, 649, 651, -1, -1, 433, 417, 653, 655, 657, 421, 423, 659, 661, 663, -1, -1, -1, -1, 665, 431, -1, -1, 435, 667, 669, 671, 673, 439, -1, -1, 443, 481, 675, 445, 447, 677, 679, 681, 683, 451, 685, 687, 689, 455, 691, 693, -1, -1, 695, 461, 697, 463, 465, 699, 701, 703, 469, 705, 707, 709, -1, -1, 711, 475, 713, 715, 717, 479, 719, 721, 483, 723, 725, 485, 727, 729, -1, -1, 731, 733, 735, 737, 739, 741, -1, -1, -1, -1, -1, -1, -1, -1, 743, 745, 747, 749, -1, -1, 751, 753, 755, 757, -1, -1, -1, -1, -1, -1, -1, -1, 759, 761, -1, -1, -1, -1, 763, 765, -1, -1, -1, -1, 767, 769, 771, 773, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 775, 777, -1, -1, -1, -1, 779, 781, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 783, 785, -1, -1, -1, -1, 787, 789, 791, 793, -1, -1, -1, -1, -1, -1, 795, 797, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 799, 801, 803, 805, -1, -1, -1, -1, 807, 809, 811, 813, -1, -1, -1, -1, 815, 817, 819, 821, -1, -1, -1, -1, 823, 825, -1, -1, 827, 829, -1, -1, -1, -1, 831, 833, -1, -1, 835, 837, 839, 841, -1, -1, -1, -1, 843, 845, 847, 849, 851, 853, 855, 857, -1, -1, -1, -1, -1, -1, 859, 861, -1, -1, -1, -1, -1, -1, 863, 865, 867, 869, -1, -1, -1, -1, 871, 873, -1, -1, -1, -1, 875, 877, -1, -1, -1, -1, 879, 881, 883, 885, 887, 889, -1, -1, -1, -1, 891, 893, -1, -1, -1, -1, 895, 897, -1, -1, -1, -1, 899, 901, 903, 905, 907, 909, 911, 913, 915, 917, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 919, 921, 923, 925, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 927, 929, 931, 933, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 935, 937, 939, 941, -1, -1, -1, -1, -1, -1, -1, -1, 943, 945, 947, 949, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 951, 953, 955, 957, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 959, 961, 963, 965, -1, -1, -1, -1, -1, -1, -1, -1, 967, 969, 971, 973, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 975, 977, 979, 981, 983, 985, 987, 989, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 991, 993, 995, 997, -1, -1, -1, -1, -1, -1, -1, -1, 999, 1001, 1003, 1005, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, 13, 15, 17, 19, 11, 21, 23, 25, 27, 29, 31, 33, 35, 37, 39, 41, 43, 45, 47, 49, 51, 53, 55, 57, 59, 61, 63, 65, 67, 69, 71, 73, 75, 77, 79, 81, 83, 85, 87, 89, 91, 93, 95, 97, 99, 101, 103, 105, 107, 109, 111, 113, 115, 117, 119, 121, 123, 125, 127, 129, 131, 133, 135, 137, 139, 141, 143, 145, 147, 149, 151, 153, 155, 157, 159, 161, 163, 165, 167, 169, 171, 173, 175, 177, 179, 181, 183, 185, 187, 189, 191, 193, 195, 197, 199, 201, 203, 205, 207, 209, 211, 213, 215, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 237, 239, 241, 243, 245, 247, 249, 251, 253, 255, 257, 259, 261, 263, 265, 267, 269, 271, 273, 275, 277, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 317, 319, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 341, 343, 345, 347, 349, 351, 353, 355, 357, 359, 361, 363, 365, 367, 369, 371, 373, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 415, 417, 419, 421, 423, 425, 427, 429, 431, 433, 435, 437, 439, 441, 443, 445, 447, 449, 451, 453, 455, 457, 459, 461, 463, 465, 467, 469, 471, 473, 475, 477, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 503, 505, 507, 509, 511, 513, 515, 517, 519, 521, 523, 525, 527, 529, 531, 533, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 555, 557, 559, 561, 563, 565, 567, 569, 571, 573, 575, 577, 579, 581, 583, 585, 587, 589, 591, 593, 595, 597, 599, 601, 603, 605, 607, 609, 611, 613, 615, 617, 619, 621, 623, 625, 627, 629, 631, 633, 635, 637, 639, 641, 643, 645, 647, 649, 651, 653, 655, 657, 659, 661, 663, 665, 667, 669, 671, 673, 675, 677, 679, 681, 683, 685, 687, 689, 691, 693, 695, 697, 699, 701, 703, 705, 707, 709, 711, 713, 715, 717, 719, 721, 723, 725, 727, 729, 731, 733, 735, 737, 739, 741, 743, 745, 747, 749, 751, 753, 755, 757, 759, 761, 763, 765, 767, 769, 771, 773, 775, 777, 779, 781, 783, 785, 787, 789, 791, 793, 795, 797, 799, 801, 803, 805, 807, 809, 811, 813, 815, 817, 819, 821, 823, 825, 827, 829, 831, 833, 835, 837, 839, 841, 843, 845, 847, 849, 851, 853, 855, 857, 859, 861, 863, 865, 867, 869, 871, 873, 875, 877, 879, 881, 883, 885, 887, 889, 891, 893, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 895, 897, 899, 901, 903, 905, 907, 909, 911, 913, 915, 917, 919, 921, 923, 925, 927, 929, 931, 933, 935, 937, 939, 941, 943, 945, 947, 949, 951, 953, 955, 957, 959, 961, 963, 965, 967, 969, 971, 973, 975, 977, 979, 981, 983, 985, 987, 989, 991, 993, 995, 997, 999, 1001, 1003, 1005, 1007, 1009, 1011, 1013, 1015, 1017, 1019, 1021, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 8, 6, 14, 12, 26, 10, 36, 22, 20, 18, 68, 84, 16, 32, 46, 58, 90, 146, 30, 114, 24, 44, 52, 190, 28, 62, 64, 42, 56, 34, 154, 140, 98, 38, 270, 134, 40, 74, 102, 108, 124, 240, 72, 48, 446, 338, 50, 176, 110, 54, 402, 168, 204, 370, 66, 60, 448, 450, 452, 198, 94, 80, 262, 164, 302, 70, 366, 414, 128, 122, 180, 76, 214, 232, 78, 152, 246, 210, 82, 188, 330, 86, 250, 318, 88, 132, 228, 92, 170, 226, 454, 96, 120, 208, 298, 326, 100, 256, 456, 104, 458, 106, 288, 202, 460, 166, 236, 292, 112, -1, -1, 384, 116, 118, 184, 304, 306, 462, 464, 382, 466, 468, 126, 470, 144, 130, 472, 196, 474, 160, 182, 350, 136, 138, 348, 310, 220, 142, 476, 478, 344, -1, -1, 148, 410, 284, 150, 322, 314, -1, -1, 156, 398, 158, 480, 308, 258, 162, 392, -1, -1, 300, 222, 212, 248, 174, 482, 362, 172, 484, 358, -1, -1, 178, 486, -1, -1, 268, 488, 490, 492, 186, 494, 224, 296, -1, -1, 192, 418, 496, 194, 316, 346, -1, -1, 498, 200, 500, 312, -1, -1, 502, 206, -1, -1, -1, -1, 504, 260, -1, -1, 394, 216, 506, 218, -1, -1, 508, 510, -1, -1, -1, -1, 512, 514, 516, 230, 518, 520, 234, 522, -1, -1, 238, 524, -1, -1, 526, 242, 528, 244, -1, -1, -1, -1, -1, -1, 252, 432, 424, 254, 530, 280, -1, -1, -1, -1, -1, -1, 264, 428, 266, 294, -1, -1, -1, -1, 272, 440, 374, 274, 276, 332, 532, 278, 534, 536, 282, 538, -1, -1, 540, 286, 542, 544, 546, 290, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 548, 550, 552, 554, 324, 556, -1, -1, 558, 560, -1, -1, 562, 564, 566, 568, 570, 320, 572, 360, 574, 576, -1, -1, 578, 328, -1, -1, -1, -1, 334, 580, 336, 582, -1, -1, 584, 340, 586, 342, -1, -1, -1, -1, 588, 590, 592, 594, 596, 352, 354, 598, 356, 600, -1, -1, -1, -1, 602, 604, 606, 364, -1, -1, 608, 368, 610, 612, 614, 372, 616, 618, 620, 376, 378, 622, 380, 624, -1, -1, -1, -1, 626, 386, 388, 628, 390, 630, -1, -1, -1, -1, 396, 632, -1, -1, 400, 634, 636, 638, 406, 404, 640, 642, 408, 644, -1, -1, 646, 412, 648, 650, 652, 416, 654, 656, 420, 658, 660, 422, 662, 664, 666, 426, 668, 670, 430, 672, -1, -1, 674, 434, 676, 436, 438, 678, -1, -1, 680, 442, 444, 682, 684, 686, 688, 690, 692, 694, 696, 698, 700, 702, 704, 706, -1, -1, 708, 710, -1, -1, -1, -1, -1, -1, -1, -1, 712, 714, -1, -1, 716, 718, -1, -1, 720, 722, -1, -1, 724, 726, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 728, 730, 732, 734, 736, 738, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 740, 742, -1, -1, -1, -1, -1, -1, -1, -1, 744, 746, -1, -1, 748, 750, 752, 754, -1, -1, -1, -1, -1, -1, 756, 758, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 760, 762, 764, 766, -1, -1, -1, -1, -1, -1, 768, 770, -1, -1, 772, 774, -1, -1, -1, -1, -1, -1, 776, 778, 780, 782, 784, 786, 788, 790, -1, -1, -1, -1, -1, -1, -1, -1, 792, 794, 796, 798, 800, 802, 804, 806, -1, -1, -1, -1, 808, 810, 812, 814, -1, -1, 816, 818, 820, 822, -1, -1, -1, -1, 824, 826, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 828, 830, 832, 834, 836, 838, 840, 842, -1, -1, -1, -1, 844, 846, 848, 850, -1, -1, -1, -1, 852, 854, -1, -1, -1, -1, -1, -1, 856, 858, 860, 862, -1, -1, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, 888, 890, 892, 894, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 896, 898, 900, 902, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 904, 906, 908, 910, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, -1, -1, -1, -1, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, -1, -1, -1, -1, 952, 954, 956, 958, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 960, 962, 964, 966, -1, -1, -1, -1, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 8, 6, 12, 18, 22, 10, 34, 50, 16, 40, 14, 46, 26, 54, 30, 20, 66, 70, 86, 24, 260, 152, 64, 98, 28, 62, 102, 254, 32, 74, 150, 36, 236, 128, 38, 114, 276, 42, 188, 108, 44, 76, 144, 48, 182, 272, 78, 460, 52, 60, 176, 56, 162, 82, 58, 328, 286, 354, 198, 118, 224, 158, 80, 416, 68, 90, 216, 72, 206, 490, 232, 324, 122, 202, 136, 492, 106, 84, 494, 294, 94, 496, 414, 348, 88, 270, 282, 92, 338, 342, 134, 96, 350, -1, -1, 100, 318, 194, 138, 244, 104, 140, 378, 498, 222, 468, 110, 430, 112, 126, 500, 116, 210, 252, 228, 120, 180, -1, -1, 124, 502, -1, -1, -1, -1, 478, 130, 132, 504, 304, 506, -1, -1, 302, 142, 508, 290, -1, -1, -1, -1, 146, 306, 148, 230, -1, -1, 172, 510, 384, 154, 156, 512, 514, 516, 364, 160, 242, 374, 450, 164, 166, 170, 168, 458, -1, -1, 518, 298, 174, 520, -1, -1, 178, 522, 248, 332, -1, -1, 390, 184, 186, 352, 346, 524, 400, 190, 192, 394, 314, 310, 526, 196, -1, -1, 200, 528, 530, 376, 204, 532, -1, -1, 534, 208, 372, 356, 536, 212, 538, 214, -1, -1, 218, 368, 268, 220, -1, -1, -1, -1, 540, 226, -1, -1, 542, 544, -1, -1, 546, 234, -1, -1, 238, 442, 420, 240, 292, 548, -1, -1, 246, 340, -1, -1, 250, 300, -1, -1, 550, 552, 454, 256, 258, 554, 556, 558, 360, 262, 264, 410, 358, 266, 560, 562, -1, -1, 564, 566, 274, 568, 570, 572, 278, 574, 280, 576, 578, 344, 284, 580, -1, -1, 288, 582, -1, -1, -1, -1, 334, 584, 428, 296, -1, -1, -1, -1, -1, -1, -1, -1, 586, 488, 588, 308, -1, -1, 312, 590, -1, -1, 316, 592, -1, -1, 320, 380, 426, 322, -1, -1, 326, 594, -1, -1, 330, 596, -1, -1, 598, 600, 602, 336, -1, -1, 604, 606, -1, -1, -1, -1, -1, -1, -1, -1, 608, 610, -1, -1, 612, 614, 616, 618, -1, -1, 620, 622, 362, 474, 624, 626, 366, 628, -1, -1, 630, 370, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 472, 382, -1, -1, 632, 386, 388, 634, -1, -1, 392, 636, 638, 640, 642, 396, 644, 398, -1, -1, 402, 646, 438, 404, 406, 408, -1, -1, -1, -1, 412, 648, 650, 652, -1, -1, 434, 418, 654, 656, 658, 422, 424, 660, 662, 664, -1, -1, -1, -1, 666, 432, -1, -1, 436, 668, 670, 672, 674, 440, -1, -1, 444, 482, 676, 446, 448, 678, 680, 682, 684, 452, 686, 688, 690, 456, 692, 694, -1, -1, 696, 462, 698, 464, 466, 700, 702, 704, 470, 706, 708, 710, -1, -1, 712, 476, 714, 716, 718, 480, 720, 722, 484, 724, 726, 486, 728, 730, -1, -1, 732, 734, 736, 738, 740, 742, -1, -1, -1, -1, -1, -1, -1, -1, 744, 746, 748, 750, -1, -1, 752, 754, 756, 758, -1, -1, -1, -1, -1, -1, -1, -1, 760, 762, -1, -1, -1, -1, 764, 766, -1, -1, -1, -1, 768, 770, 772, 774, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 776, 778, -1, -1, -1, -1, 780, 782, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 784, 786, -1, -1, -1, -1, 788, 790, 792, 794, -1, -1, -1, -1, -1, -1, 796, 798, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 800, 802, 804, 806, -1, -1, -1, -1, 808, 810, 812, 814, -1, -1, -1, -1, 816, 818, 820, 822, -1, -1, -1, -1, 824, 826, -1, -1, 828, 830, -1, -1, -1, -1, 832, 834, -1, -1, 836, 838, 840, 842, -1, -1, -1, -1, 844, 846, 848, 850, 852, 854, 856, 858, -1, -1, -1, -1, -1, -1, 860, 862, -1, -1, -1, -1, -1, -1, 864, 866, 868, 870, -1, -1, -1, -1, 872, 874, -1, -1, -1, -1, 876, 878, -1, -1, -1, -1, 880, 882, 884, 886, 888, 890, -1, -1, -1, -1, 892, 894, -1, -1, -1, -1, 896, 898, -1, -1, -1, -1, 900, 902, 904, 906, 908, 910, 912, 914, 916, 918, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 920, 922, 924, 926, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 928, 930, 932, 934, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 936, 938, 940, 942, -1, -1, -1, -1, -1, -1, -1, -1, 944, 946, 948, 950, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 952, 954, 956, 958, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 960, 962, 964, 966, -1, -1, -1, -1, -1, -1, -1, -1, 968, 970, 972, 974, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 976, 978, 980, 982, 984, 986, 988, 990, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 992, 994, 996, 998, -1, -1, -1, -1, -1, -1, -1, -1, 1000, 1002, 1004, 1006, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, 14, 16, 18, 20, 12, 22, 24, 26, 28, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90, 92, 94, 96, 98, 100, 102, 104, 106, 108, 110, 112, 114, 116, 118, 120, 122, 124, 126, 128, 130, 132, 134, 136, 138, 140, 142, 144, 146, 148, 150, 152, 154, 156, 158, 160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 180, 182, 184, 186, 188, 190, 192, 194, 196, 198, 200, 202, 204, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, 432, 434, 436, 438, 440, 442, 444, 446, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, 512, 514, 516, 518, 520, 522, 524, 526, 528, 530, 532, 534, 536, 538, 540, 542, 544, 546, 548, 550, 552, 554, 556, 558, 560, 562, 564, 566, 568, 570, 572, 574, 576, 578, 580, 582, 584, 586, 588, 590, 592, 594, 596, 598, 600, 602, 604, 606, 608, 610, 612, 614, 616, 618, 620, 622, 624, 626, 628, 630, 632, 634, 636, 638, 640, 642, 644, 646, 648, 650, 652, 654, 656, 658, 660, 662, 664, 666, 668, 670, 672, 674, 676, 678, 680, 682, 684, 686, 688, 690, 692, 694, 696, 698, 700, 702, 704, 706, 708, 710, 712, 714, 716, 718, 720, 722, 724, 726, 728, 730, 732, 734, 736, 738, 740, 742, 744, 746, 748, 750, 752, 754, 756, 758, 760, 762, 764, 766, 768, 770, 772, 774, 776, 778, 780, 782, 784, 786, 788, 790, 792, 794, 796, 798, 800, 802, 804, 806, 808, 810, 812, 814, 816, 818, 820, 822, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 850, 852, 854, 856, 858, 860, 862, 864, 866, 868, 870, 872, 874, 876, 878, 880, 882, 884, 886, 888, 890, 892, 894, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 896, 898, 900, 902, 904, 906, 908, 910, 912, 914, 916, 918, 920, 922, 924, 926, 928, 930, 932, 934, 936, 938, 940, 942, 944, 946, 948, 950, 952, 954, 956, 958, 960, 962, 964, 966, 968, 970, 972, 974, 976, 978, 980, 982, 984, 986, 988, 990, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 5, 5, 4, 4, 14, 14, 11, 11, 10, 10, 9, 9, 22, 22, 6, 6, 26, 26, 20, 20, 15, 15, 31, 31, 8, 8, 35, 35, 38, 38, 29, 29, 23, 23, 16, 16, 45, 45, 48, 48, 24, 24, 51, 51, 30, 30, 17, 17, 57, 57, 27, 27, 28, 28, 56, 56, 12, 12, 67, 67, 44, 44, 39, 39, 73, 73, 76, 76, 63, 63, 80, 80, 13, 13, 83, 83, 86, 86, 18, 18, 89, 89, 62, 62, 93, 93, 34, 34, 98, 98, 40, 40, 101, 101, 103, 103, 41, 41, 50, 50, 110, 110, 21, 21, 114, 114, 115, 115, 94, 94, 71, 71, 42, 42, 124, 124, 70, 70, 127, 127, 87, 87, 37, 37, 134, 134, 135, 135, 33, 33, 139, 139, 126, 126, 19, 19, 145, 145, 148, 148, 77, 77, 32, 32, 153, 153, 155, 155, 131, 131, 159, 159, 65, 65, 107, 107, 53, 53, 90, 90, 170, 170, 167, 167, 49, 49, 175, 175, 72, 72, 132, 132, 116, 116, 183, 183, 81, 81, 25, 25, 189, 189, 192, 192, 129, 129, 61, 61, 198, 198, 105, 105, 54, 54, 204, 204, 95, 95, 79, 79, 165, 165, 74, 74, 214, 214, 216, 216, 138, 138, 164, 164, 185, 185, 91, 91, 88, 88, 228, 228, 75, 75, 231, 231, 108, 108, 235, 235, 43, 43, 240, 240, 242, 242, 78, 78, 166, 166, 84, 84, 249, 249, 252, 252, 99, 99, 158, 158, 210, 210, 64, 64, 261, 261, 263, 263, 179, 179, 36, 36, 269, 269, 272, 272, 273, 273, 276, 276, 254, 254, 279, 279, 147, 147, 284, 284, 104, 104, 288, 288, 109, 109, 264, 264, 186, 186, 96, 96, 163, 163, 66, 66, 117, 117, 118, 118, 157, 157, 137, 137, 200, 200, 150, 150, 193, 193, 85, 85, 318, 318, 149, 149, 305, 305, 97, 97, 326, 326, 82, 82, 274, 274, 331, 331, 333, 333, 47, 47, 338, 338, 340, 340, 142, 142, 194, 194, 136, 136, 133, 133, 350, 350, 351, 351, 353, 353, 172, 172, 320, 320, 169, 169, 362, 362, 68, 68, 366, 366, 55, 55, 370, 370, 271, 271, 374, 374, 375, 375, 377, 377, 121, 121, 113, 113, 384, 384, 385, 385, 387, 387, 160, 160, 213, 213, 393, 393, 154, 154, 397, 397, 52, 52, 402, 402, 401, 401, 405, 405, 146, 146, 410, 410, 69, 69, 414, 414, 190, 190, 417, 417, 420, 420, 251, 251, 424, 424, 262, 262, 427, 427, 250, 250, 432, 432, 434, 434, 435, 435, 270, 270, 440, 440, 441, 441, 46, 46, 58, 58, 59, 59, 60, 60, 92, 92, 100, 100, 102, 102, 106, 106, 119, 119, 120, 120, 122, 122, 123, 123, 125, 125, 128, 128, 130, 130, 140, 140, 141, 141, 156, 156, 168, 168, 171, 171, 176, 176, 180, 180, 181, 181, 182, 182, 184, 184, 191, 191, 197, 197, 199, 199, 203, 203, 209, 209, 215, 215, 219, 219, 220, 220, 225, 225, 226, 226, 227, 227, 229, 229, 230, 230, 232, 232, 236, 236, 239, 239, 241, 241, 253, 253, 275, 275, 277, 277, 278, 278, 280, 280, 283, 283, 285, 285, 286, 286, 287, 287, 301, 301, 302, 302, 303, 303, 304, 304, 306, 306, 309, 309, 310, 310, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 319, 319, 321, 321, 322, 322, 325, 325, 332, 332, 334, 334, 337, 337, 339, 339, 345, 345, 346, 346, 347, 347, 348, 348, 349, 349, 352, 352, 354, 354, 359, 359, 360, 360, 361, 361, 365, 365, 367, 367, 368, 368, 369, 369, 371, 371, 372, 372, 373, 373, 376, 376, 378, 378, 383, 383, 386, 386, 388, 388, 394, 394, 398, 398, 399, 399, 400, 400, 403, 403, 404, 404, 406, 406, 409, 409, 411, 411, 412, 412, 413, 413, 415, 415, 416, 416, 418, 418, 419, 419, 421, 421, 422, 422, 423, 423, 425, 425, 426, 426, 428, 428, 431, 431, 433, 433, 436, 436, 439, 439, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446, 447, 447, 448, 448, 449, 449, 450, 450, 451, 451, 452, 452, 453, 453, 454, 454, 457, 457, 458, 458, 467, 467, 468, 468, 471, 471, 472, 472, 475, 475, 476, 476, 479, 479, 480, 480, 493, 493, 494, 494, 495, 495, 496, 496, 497, 497, 498, 498, 515, 515, 516, 516, 525, 525, 526, 526, 529, 529, 530, 530, 531, 531, 532, 532, 539, 539, 540, 540, 569, 569, 570, 570, 571, 571, 572, 572, 579, 579, 580, 580, 583, 583, 584, 584, 591, 591, 592, 592, 593, 593, 594, 594, 595, 595, 596, 596, 597, 597, 598, 598, 607, 607, 608, 608, 609, 609, 610, 610, 611, 611, 612, 612, 613, 613, 614, 614, 619, 619, 620, 620, 621, 621, 622, 622, 625, 625, 626, 626, 627, 627, 628, 628, 633, 633, 634, 634, 645, 645, 646, 646, 647, 647, 648, 648, 649, 649, 650, 650, 651, 651, 652, 652, 657, 657, 658, 658, 659, 659, 660, 660, 665, 665, 666, 666, 673, 673, 674, 674, 675, 675, 676, 676, 679, 679, 680, 680, 681, 681, 682, 682, 683, 683, 684, 684, 685, 685, 686, 686, 687, 687, 688, 688, 689, 689, 690, 690, 691, 691, 692, 692, 693, 693, 694, 694, 707, 707, 708, 708, 709, 709, 710, 710, 731, 731, 732, 732, 733, 733, 734, 734, 759, 759, 760, 760, 761, 761, 762, 762, 783, 783, 784, 784, 785, 785, 786, 786, 791, 791, 792, 792, 793, 793, 794, 794, 807, 807, 808, 808, 809, 809, 810, 810, 815, 815, 816, 816, 817, 817, 818, 818, 827, 827, 828, 828, 829, 829, 830, 830, 843, 843, 844, 844, 845, 845, 846, 846, 855, 855, 856, 856, 857, 857, 858, 858, 863, 863, 864, 864, 865, 865, 866, 866, 867, 867, 868, 868, 869, 869, 870, 870, 879, 879, 880, 880, 881, 881, 882, 882, 883, 883, 884, 884, 885, 885, 886, 886, 975, 975, 976, 976, 977, 977, 978, 978, 979, 979, 980, 980, 981, 981, 982, 982),
                (-1, 0, 0, 1, 1, 3, 3, 2, 2, 7, 7, 4, 4, 12, 12, 10, 10, 5, 5, 17, 17, 6, 6, 21, 21, 14, 14, 26, 26, 16, 16, 30, 30, 8, 8, 33, 33, 36, 36, 11, 11, 39, 39, 42, 42, 13, 13, 45, 45, 9, 9, 50, 50, 15, 15, 53, 53, 56, 56, 51, 51, 27, 27, 24, 24, 18, 18, 66, 66, 19, 19, 69, 69, 31, 31, 43, 43, 48, 48, 64, 64, 55, 55, 79, 79, 20, 20, 86, 86, 67, 67, 89, 89, 82, 82, 93, 93, 25, 25, 97, 97, 28, 28, 102, 102, 78, 78, 41, 41, 108, 108, 110, 110, 37, 37, 113, 113, 61, 61, 117, 117, 74, 74, 121, 121, 111, 111, 35, 35, 128, 128, 129, 129, 92, 92, 76, 76, 100, 100, 103, 103, 136, 136, 44, 44, 143, 143, 145, 145, 32, 32, 23, 23, 152, 152, 153, 153, 63, 63, 158, 158, 54, 54, 162, 162, 163, 163, 165, 165, 164, 164, 149, 149, 171, 171, 52, 52, 175, 175, 118, 118, 46, 46, 182, 182, 183, 183, 40, 40, 188, 188, 189, 189, 99, 99, 194, 194, 60, 60, 197, 197, 75, 75, 201, 201, 70, 70, 206, 206, 114, 114, 210, 210, 212, 212, 68, 68, 215, 215, 218, 218, 106, 106, 62, 62, 224, 224, 116, 116, 146, 146, 72, 72, 232, 232, 34, 34, 235, 235, 238, 238, 159, 159, 101, 101, 243, 243, 177, 177, 247, 247, 115, 115, 29, 29, 254, 254, 255, 255, 22, 22, 260, 260, 261, 261, 264, 264, 217, 217, 87, 87, 47, 47, 271, 271, 38, 38, 275, 275, 277, 277, 88, 88, 281, 281, 58, 58, 285, 285, 138, 138, 239, 239, 81, 81, 294, 294, 170, 170, 248, 248, 135, 135, 131, 131, 144, 144, 306, 306, 192, 192, 309, 309, 191, 191, 313, 313, 98, 98, 317, 317, 320, 320, 73, 73, 323, 323, 57, 57, 327, 327, 178, 178, 291, 291, 334, 334, 90, 90, 244, 244, 91, 91, 280, 280, 185, 185, 85, 85, 94, 94, 184, 184, 59, 59, 208, 208, 263, 263, 259, 259, 359, 359, 157, 157, 363, 363, 216, 216, 368, 368, 207, 207, 160, 160, 200, 200, 104, 104, 318, 318, 380, 380, 151, 151, 384, 384, 385, 385, 181, 181, 389, 389, 190, 190, 394, 394, 396, 396, 187, 187, 399, 399, 402, 402, 403, 403, 404, 404, 262, 262, 409, 409, 84, 84, 65, 65, 416, 416, 237, 237, 420, 420, 421, 421, 319, 319, 293, 293, 109, 109, 430, 430, 415, 415, 433, 433, 401, 401, 438, 438, 236, 236, 441, 441, 444, 444, 445, 445, 161, 161, 450, 450, 253, 253, 454, 454, 166, 166, 49, 49, 460, 460, 462, 462, 463, 463, 107, 107, 467, 467, 379, 379, 360, 360, 474, 474, 127, 127, 478, 478, 442, 442, 481, 481, 484, 484, 304, 304, 71, 71, 77, 77, 80, 80, 83, 83, 105, 105, 112, 112, 122, 122, 130, 130, 132, 132, 137, 137, 150, 150, 154, 154, 155, 155, 156, 156, 169, 169, 172, 172, 176, 176, 186, 186, 193, 193, 198, 198, 199, 199, 202, 202, 205, 205, 209, 209, 211, 211, 223, 223, 227, 227, 228, 228, 231, 231, 240, 240, 251, 251, 252, 252, 256, 256, 257, 257, 258, 258, 265, 265, 266, 266, 269, 269, 270, 270, 272, 272, 273, 273, 274, 274, 276, 276, 278, 278, 279, 279, 282, 282, 286, 286, 292, 292, 303, 303, 305, 305, 310, 310, 314, 314, 324, 324, 328, 328, 331, 331, 332, 332, 333, 333, 337, 337, 338, 338, 347, 347, 348, 348, 351, 351, 352, 352, 353, 353, 354, 354, 357, 357, 358, 358, 361, 361, 362, 362, 364, 364, 367, 367, 383, 383, 386, 386, 390, 390, 391, 391, 392, 392, 393, 393, 395, 395, 400, 400, 410, 410, 411, 411, 412, 412, 417, 417, 418, 418, 419, 419, 422, 422, 423, 423, 424, 424, 429, 429, 434, 434, 435, 435, 436, 436, 437, 437, 443, 443, 446, 446, 447, 447, 448, 448, 449, 449, 451, 451, 452, 452, 453, 453, 455, 455, 456, 456, 459, 459, 461, 461, 464, 464, 465, 465, 466, 466, 468, 468, 469, 469, 470, 470, 473, 473, 475, 475, 476, 476, 477, 477, 479, 479, 480, 480, 482, 482, 483, 483, 485, 485, 486, 486, 489, 489, 490, 490, 491, 491, 492, 492, 493, 493, 494, 494, 503, 503, 504, 504, 505, 505, 506, 506, 509, 509, 510, 510, 511, 511, 512, 512, 521, 521, 522, 522, 527, 527, 528, 528, 533, 533, 534, 534, 535, 535, 536, 536, 547, 547, 548, 548, 553, 553, 554, 554, 567, 567, 568, 568, 573, 573, 574, 574, 575, 575, 576, 576, 583, 583, 584, 584, 607, 607, 608, 608, 609, 609, 610, 610, 615, 615, 616, 616, 617, 617, 618, 618, 623, 623, 624, 624, 625, 625, 626, 626, 631, 631, 632, 632, 635, 635, 636, 636, 641, 641, 642, 642, 645, 645, 646, 646, 647, 647, 648, 648, 653, 653, 654, 654, 655, 655, 656, 656, 657, 657, 658, 658, 659, 659, 660, 660, 667, 667, 668, 668, 675, 675, 676, 676, 677, 677, 678, 678, 683, 683, 684, 684, 689, 689, 690, 690, 695, 695, 696, 696, 697, 697, 698, 698, 699, 699, 700, 700, 705, 705, 706, 706, 711, 711, 712, 712, 717, 717, 718, 718, 719, 719, 720, 720, 721, 721, 722, 722, 723, 723, 724, 724, 725, 725, 726, 726, 743, 743, 744, 744, 745, 745, 746, 746, 759, 759, 760, 760, 761, 761, 762, 762, 775, 775, 776, 776, 777, 777, 778, 778, 787, 787, 788, 788, 789, 789, 790, 790, 835, 835, 836, 836, 837, 837, 838, 838, 851, 851, 852, 852, 853, 853, 854, 854, 863, 863, 864, 864, 865, 865, 866, 866, 879, 879, 880, 880, 881, 881, 882, 882, 883, 883, 884, 884, 885, 885, 886, 886, 899, 899, 900, 900, 901, 901, 902, 902, 911, 911, 912, 912, 913, 913, 914, 914, 975, 975, 976, 976, 977, 977, 978, 978, 979, 979, 980, 980, 981, 981, 982, 982),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 10, 10, 11, 11, 12, 12, 13, 13, 14, 14, 15, 15, 16, 16, 17, 17, 18, 18, 19, 19, 20, 20, 21, 21, 22, 22, 23, 23, 24, 24, 25, 25, 26, 26, 27, 27, 28, 28, 29, 29, 30, 30, 31, 31, 32, 32, 33, 33, 34, 34, 35, 35, 36, 36, 37, 37, 38, 38, 39, 39, 40, 40, 41, 41, 42, 42, 43, 43, 44, 44, 45, 45, 46, 46, 47, 47, 48, 48, 49, 49, 50, 50, 51, 51, 52, 52, 53, 53, 54, 54, 55, 55, 56, 56, 57, 57, 58, 58, 59, 59, 60, 60, 61, 61, 62, 62, 63, 63, 64, 64, 65, 65, 66, 66, 67, 67, 68, 68, 69, 69, 70, 70, 71, 71, 72, 72, 73, 73, 74, 74, 75, 75, 76, 76, 77, 77, 78, 78, 79, 79, 80, 80, 81, 81, 82, 82, 83, 83, 84, 84, 85, 85, 86, 86, 87, 87, 88, 88, 89, 89, 90, 90, 91, 91, 92, 92, 93, 93, 94, 94, 95, 95, 96, 96, 97, 97, 98, 98, 99, 99, 100, 100, 101, 101, 102, 102, 103, 103, 104, 104, 105, 105, 106, 106, 107, 107, 108, 108, 109, 109, 110, 110, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 117, 117, 118, 118, 119, 119, 120, 120, 121, 121, 122, 122, 123, 123, 124, 124, 125, 125, 126, 126, 127, 127, 128, 128, 129, 129, 130, 130, 131, 131, 132, 132, 133, 133, 134, 134, 135, 135, 136, 136, 137, 137, 138, 138, 139, 139, 140, 140, 141, 141, 142, 142, 143, 143, 144, 144, 145, 145, 146, 146, 147, 147, 148, 148, 149, 149, 150, 150, 151, 151, 152, 152, 153, 153, 154, 154, 155, 155, 156, 156, 157, 157, 158, 158, 159, 159, 160, 160, 161, 161, 162, 162, 163, 163, 164, 164, 165, 165, 166, 166, 167, 167, 168, 168, 169, 169, 170, 170, 171, 171, 172, 172, 173, 173, 174, 174, 175, 175, 176, 176, 177, 177, 178, 178, 179, 179, 180, 180, 181, 181, 182, 182, 183, 183, 184, 184, 185, 185, 186, 186, 187, 187, 188, 188, 189, 189, 190, 190, 191, 191, 192, 192, 193, 193, 194, 194, 195, 195, 196, 196, 197, 197, 198, 198, 199, 199, 200, 200, 201, 201, 202, 202, 203, 203, 204, 204, 205, 205, 206, 206, 207, 207, 208, 208, 209, 209, 210, 210, 211, 211, 212, 212, 213, 213, 214, 214, 215, 215, 216, 216, 217, 217, 218, 218, 219, 219, 220, 220, 221, 221, 222, 222, 223, 223, 224, 224, 225, 225, 226, 226, 227, 227, 228, 228, 229, 229, 230, 230, 231, 231, 232, 232, 233, 233, 234, 234, 235, 235, 236, 236, 237, 237, 238, 238, 239, 239, 240, 240, 241, 241, 242, 242, 243, 243, 244, 244, 245, 245, 246, 246, 247, 247, 248, 248, 249, 249, 250, 250, 251, 251, 252, 252, 253, 253, 254, 254, 255, 255, 256, 256, 257, 257, 258, 258, 259, 259, 260, 260, 261, 261, 262, 262, 263, 263, 264, 264, 265, 265, 266, 266, 267, 267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 272, 273, 273, 274, 274, 275, 275, 276, 276, 277, 277, 278, 278, 279, 279, 280, 280, 281, 281, 282, 282, 283, 283, 284, 284, 285, 285, 286, 286, 287, 287, 288, 288, 289, 289, 290, 290, 291, 291, 292, 292, 293, 293, 294, 294, 295, 295, 296, 296, 297, 297, 298, 298, 299, 299, 300, 300, 301, 301, 302, 302, 303, 303, 304, 304, 305, 305, 306, 306, 307, 307, 308, 308, 309, 309, 310, 310, 311, 311, 312, 312, 313, 313, 314, 314, 315, 315, 316, 316, 317, 317, 318, 318, 319, 319, 320, 320, 321, 321, 322, 322, 323, 323, 324, 324, 325, 325, 326, 326, 327, 327, 328, 328, 329, 329, 330, 330, 331, 331, 332, 332, 333, 333, 334, 334, 335, 335, 336, 336, 337, 337, 338, 338, 339, 339, 340, 340, 341, 341, 342, 342, 343, 343, 344, 344, 345, 345, 346, 346, 347, 347, 348, 348, 349, 349, 350, 350, 351, 351, 352, 352, 353, 353, 354, 354, 355, 355, 356, 356, 357, 357, 358, 358, 359, 359, 360, 360, 361, 361, 362, 362, 363, 363, 364, 364, 365, 365, 366, 366, 367, 367, 368, 368, 369, 369, 370, 370, 371, 371, 372, 372, 373, 373, 374, 374, 375, 375, 376, 376, 377, 377, 378, 378, 379, 379, 380, 380, 381, 381, 382, 382, 383, 383, 384, 384, 385, 385, 386, 386, 387, 387, 388, 388, 389, 389, 390, 390, 391, 391, 392, 392, 393, 393, 394, 394, 395, 395, 396, 396, 397, 397, 398, 398, 399, 399, 400, 400, 401, 401, 402, 402, 403, 403, 404, 404, 405, 405, 406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 412, 412, 413, 413, 414, 414, 415, 415, 416, 416, 417, 417, 418, 418, 419, 419, 420, 420, 421, 421, 422, 422, 423, 423, 424, 424, 425, 425, 426, 426, 427, 427, 428, 428, 429, 429, 430, 430, 431, 431, 432, 432, 433, 433, 434, 434, 435, 435, 436, 436, 437, 437, 438, 438, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 444, 444, 445, 445, 446, 446, 703, 703, 704, 704, 705, 705, 706, 706, 707, 707, 708, 708, 709, 709, 710, 710, 711, 711, 712, 712, 713, 713, 714, 714, 715, 715, 716, 716, 717, 717, 718, 718, 719, 719, 720, 720, 721, 721, 722, 722, 723, 723, 724, 724, 725, 725, 726, 726, 727, 727, 728, 728, 729, 729, 730, 730, 731, 731, 732, 732, 733, 733, 734, 734, 735, 735, 736, 736, 737, 737, 738, 738, 739, 739, 740, 740, 741, 741, 742, 742, 743, 743, 744, 744, 745, 745, 746, 746, 747, 747, 748, 748, 749, 749, 750, 750, 751, 751, 752, 752, 753, 753, 754, 754, 755, 755, 756, 756, 757, 757, 758, 758, 759, 759, 760, 760, 761, 761, 762, 762, 763, 763, 764, 764, 765, 765, 766, 766)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 4, 4, 3, 3, 4, 4, 5, 5, 4, 4, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 5, 5, 6, 6, 3, 3, 4, 4, 5, 5, 6, 6, 6, 6, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 6, 6, 6, 6, 7, 7, 6, 6, 6, 6, 7, 7, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 4, 4, 5, 5, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 5, 5, 6, 6, 7, 7, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 4, 4, 5, 5, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 7, 7, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 8, 8, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 5, 5, 5, 5, 6, 6, 5, 5, 6, 6, 3, 3, 4, 4, 5, 5, 4, 4, 5, 5, 6, 6, 5, 5, 6, 6, 4, 4, 5, 5, 5, 5, 6, 6, 7, 7, 6, 6, 7, 7, 6, 6, 5, 5, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 6, 6, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 5, 5, 6, 6, 7, 7, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 6, 6, 7, 7, 9, 9, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 4, 4, 5, 5, 6, 6, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 6, 6, 7, 7, 8, 8, 5, 5, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 7, 7, 8, 8, 6, 6, 7, 7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 8, 8, 7, 7, 9, 9, 8, 8, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 5, 5, 6, 6, 7, 7, 8, 8, 7, 7, 8, 8, 9, 9, 7, 7, 8, 8, 6, 6, 7, 7, 6, 6, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 6, 6, 7, 7, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 7, 7, 8, 8, 8, 8, 7, 7, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((111, 112, 143, 144, 151, 152, 161, 162, 173, 174, 177, 178, 187, 188, 195, 196, 201, 202, 205, 206, 207, 208, 211, 212, 217, 218, 221, 222, 223, 224, 233, 234, 237, 238, 243, 244, 245, 246, 247, 248, 255, 256, 257, 258, 259, 260, 265, 266, 267, 268, 281, 282, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 307, 308, 311, 312, 323, 324, 327, 328, 329, 330, 335, 336, 341, 342, 343, 344, 355, 356, 357, 358, 363, 364, 379, 380, 381, 382, 389, 390, 391, 392, 395, 396, 407, 408, 429, 430, 437, 438, 455, 456, 459, 460, 461, 462, 463, 464, 465, 466, 469, 470, 473, 474, 477, 478, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 517, 518, 519, 520, 521, 522, 523, 524, 527, 528, 533, 534, 535, 536, 537, 538, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 573, 574, 575, 576, 577, 578, 581, 582, 585, 586, 587, 588, 589, 590, 599, 600, 601, 602, 603, 604, 605, 606, 615, 616, 617, 618, 623, 624, 629, 630, 631, 632, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 653, 654, 655, 656, 661, 662, 663, 664, 667, 668, 669, 670, 671, 672, 677, 678, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 763, 764, 765, 766, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 787, 788, 789, 790, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 811, 812, 813, 814, 819, 820, 821, 822, 823, 824, 825, 826, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 847, 848, 849, 850, 851, 852, 853, 854, 859, 860, 861, 862, 871, 872, 873, 874, 875, 876, 877, 878, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (95, 96, 119, 120, 123, 124, 125, 126, 133, 134, 139, 140, 141, 142, 147, 148, 167, 168, 173, 174, 179, 180, 195, 196, 203, 204, 213, 214, 219, 220, 221, 222, 225, 226, 229, 230, 233, 234, 241, 242, 245, 246, 249, 250, 267, 268, 283, 284, 287, 288, 289, 290, 295, 296, 297, 298, 299, 300, 301, 302, 307, 308, 311, 312, 315, 316, 321, 322, 325, 326, 329, 330, 335, 336, 339, 340, 341, 342, 343, 344, 345, 346, 349, 350, 355, 356, 365, 366, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 381, 382, 387, 388, 397, 398, 405, 406, 407, 408, 413, 414, 425, 426, 427, 428, 431, 432, 439, 440, 457, 458, 471, 472, 487, 488, 495, 496, 497, 498, 499, 500, 501, 502, 507, 508, 513, 514, 515, 516, 517, 518, 519, 520, 523, 524, 525, 526, 529, 530, 531, 532, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 549, 550, 551, 552, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 569, 570, 571, 572, 577, 578, 579, 580, 581, 582, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 611, 612, 613, 614, 619, 620, 621, 622, 627, 628, 629, 630, 633, 634, 637, 638, 639, 640, 643, 644, 649, 650, 651, 652, 661, 662, 663, 664, 665, 666, 669, 670, 671, 672, 673, 674, 679, 680, 681, 682, 685, 686, 687, 688, 691, 692, 693, 694, 701, 702, 703, 704, 707, 708, 709, 710, 713, 714, 715, 716, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 763, 764, 765, 766, 767, 768, 769, 770, 771, 772, 773, 774, 779, 780, 781, 782, 783, 784, 785, 786, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 855, 856, 857, 858, 859, 860, 861, 862, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 903, 904, 905, 906, 907, 908, 909, 910, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022),
                (447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 767, 768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 863, 864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 2, 1, 0, -2, -2, 1, -2, -2, 2, 0, -2, -2, 0, -2, -2, 1, 0, 2, -2, -2, 1, -2, -2, 2, 1, -2, -2, 0, -2, -2, 2, 2, 0, 1, -2, -2, 1, -2, -2, 0, 1, -2, -2, 1, -2, -2, 0, 1, 2, -2, -2, 0, -2, -2, 1, 2, -2, -2, 0, -2, -2),
                (1, 0, 1, 0, 0, -2, -2, 0, -2, -2, 0, 2, -2, -2, 2, -2, -2, 1, 0, 2, -2, -2, 2, -2, -2, 2, 1, -2, -2, 1, -2, -2, 1, 2, 0, 1, -2, -2, 1, -2, -2, 2, 2, -2, -2, 0, -2, -2, 0, 2, 2, -2, -2, 1, -2, -2, 0, 0, -2, -2, 2, -2, -2),
                (1, 0, 1, 2, 0, -2, -2, 2, -2, -2, 1, 2, -2, -2, 1, -2, -2, 0, 1, 2, -2, -2, 2, -2, -2, 0, 1, -2, -2, 0, -2, -2, 2, 0, 2, 0, -2, -2, 0, -2, -2, 2, 1, -2, -2, 1, -2, -2, 0, 2, 1, -2, -2, 1, -2, -2, 1, 2, -2, -2, 0, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((2234, 134, 92, 1637, 13351, -256, -256, 1638, -256, -256, 109, 16424, -256, -256, 12547, -256, -256, 1558, 6389, 164, -256, -256, 1143, -256, -256, 164, 1818, -256, -256, 19242, -256, -256, 109, 92, 63846, 2595, -256, -256, 3072, -256, -256, 57532, 2650, -256, -256, 3356, -256, -256, 43416, 2840, 134, -256, -256, 37491, -256, -256, 3227, 134, -256, -256, 61303, -256, -256),
                (2452, 15589, 1124, 3885, 1243, -256, -256, 10054, -256, -256, 11452, 134, -256, -256, 134, -256, -256, 1870, 22400, 92, -256, -256, 92, -256, -256, 134, 2234, -256, -256, 2364, -256, -256, 3039, 92, 53674, 2580, -256, -256, 2794, -256, -256, 134, 109, -256, -256, 33359, -256, -256, 60159, 134, 109, -256, -256, 3532, -256, -256, 75727, 68030, -256, -256, 92, -256, -256),
                (2362, 17552, 1120, 134, 3928, -256, -256, 164, -256, -256, 1438, 164, -256, -256, 1655, -256, -256, 28255, 1831, 92, -256, -256, 134, -256, -256, 35639, 2208, -256, -256, 39738, -256, -256, 134, 61177, 109, 49287, -256, -256, 47666, -256, -256, 92, 3068, -256, -256, 3369, -256, -256, 39772, 164, 2589, -256, -256, 2847, -256, -256, 3112, 164, -256, -256, 48394, -256, -256)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((38, 41, 40, 40, 41, 17, 43, 37, 0, 37, 40, 40, 15, 42, 41, 13, 42, 41, 42, 13, 12, 14, 43, 43, 42, 39, 39, 40, 39, 40, 4, 43, 34, 33, 32, 4, 13, 1, 41, 43, 40, 33, 6, 14, 1, 42, 42, 39, 36, 6, 11, 6, 14, 1, 0, 6, 42, 42, 42, 43, 41, 22, 43),
                (38, 40, 16, 30, 9, 0, 16, 39, 36, 43, 3, 0, 0, 0, 10, 5, 16, 42, 43, 39, 34, 41, 43, 43, 43, 41, 40, 41, 39, 42, 42, 40, 34, 36, 32, 1, 3, 0, 42, 43, 41, 36, 36, 35, 36, 37, 2, 42, 32, 4, 1, 0, 2, 9, 10, 3, 41, 29, 25, 33, 42, 42, 43),
                (38, 41, 18, 32, 30, 9, 39, 34, 34, 34, 4, 11, 9, 19, 2, 5, 0, 42, 35, 42, 39, 42, 12, 5, 27, 43, 41, 42, 22, 43, 42, 43, 34, 33, 5, 4, 1, 15, 8, 3, 27, 42, 41, 43, 38, 42, 43, 41, 36, 4, 3, 10, 1, 5, 13, 1, 42, 43, 43, 43, 41, 13, 43)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 2, 3, 4, 5, -1, -1, 8, -1, -1, 11, 12, -1, -1, 15, -1, -1, 18, 19, 20, -1, -1, 23, -1, -1, 26, 27, -1, -1, 30, -1, -1, 33, 34, 35, 36, -1, -1, 39, -1, -1, 42, 43, -1, -1, 46, -1, -1, 49, 50, 51, -1, -1, 54, -1, -1, 57, 58, -1, -1, 61, -1, -1),
                (1, 2, 3, 4, 5, -1, -1, 8, -1, -1, 11, 12, -1, -1, 15, -1, -1, 18, 19, 20, -1, -1, 23, -1, -1, 26, 27, -1, -1, 30, -1, -1, 33, 34, 35, 36, -1, -1, 39, -1, -1, 42, 43, -1, -1, 46, -1, -1, 49, 50, 51, -1, -1, 54, -1, -1, 57, 58, -1, -1, 61, -1, -1),
                (1, 2, 3, 4, 5, -1, -1, 8, -1, -1, 11, 12, -1, -1, 15, -1, -1, 18, 19, 20, -1, -1, 23, -1, -1, 26, 27, -1, -1, 30, -1, -1, 33, 34, 35, 36, -1, -1, 39, -1, -1, 42, 43, -1, -1, 46, -1, -1, 49, 50, 51, -1, -1, 54, -1, -1, 57, 58, -1, -1, 61, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((32, 17, 10, 7, 6, -1, -1, 9, -1, -1, 14, 13, -1, -1, 16, -1, -1, 25, 22, 21, -1, -1, 24, -1, -1, 29, 28, -1, -1, 31, -1, -1, 48, 41, 38, 37, -1, -1, 40, -1, -1, 45, 44, -1, -1, 47, -1, -1, 56, 53, 52, -1, -1, 55, -1, -1, 60, 59, -1, -1, 62, -1, -1),
                (32, 17, 10, 7, 6, -1, -1, 9, -1, -1, 14, 13, -1, -1, 16, -1, -1, 25, 22, 21, -1, -1, 24, -1, -1, 29, 28, -1, -1, 31, -1, -1, 48, 41, 38, 37, -1, -1, 40, -1, -1, 45, 44, -1, -1, 47, -1, -1, 56, 53, 52, -1, -1, 55, -1, -1, 60, 59, -1, -1, 62, -1, -1),
                (32, 17, 10, 7, 6, -1, -1, 9, -1, -1, 14, 13, -1, -1, 16, -1, -1, 25, 22, 21, -1, -1, 24, -1, -1, 29, 28, -1, -1, 31, -1, -1, 48, 41, 38, 37, -1, -1, 40, -1, -1, 45, 44, -1, -1, 47, -1, -1, 56, 53, 52, -1, -1, 55, -1, -1, 60, 59, -1, -1, 62, -1, -1)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 1, 2, 3, 4, 4, 3, 7, 7, 2, 10, 11, 11, 10, 14, 14, 1, 17, 18, 19, 19, 18, 22, 22, 17, 25, 26, 26, 25, 29, 29, 0, 32, 33, 34, 35, 35, 34, 38, 38, 33, 41, 42, 42, 41, 45, 45, 32, 48, 49, 50, 50, 49, 53, 53, 48, 56, 57, 57, 56, 60, 60),
                (-1, 0, 1, 2, 3, 4, 4, 3, 7, 7, 2, 10, 11, 11, 10, 14, 14, 1, 17, 18, 19, 19, 18, 22, 22, 17, 25, 26, 26, 25, 29, 29, 0, 32, 33, 34, 35, 35, 34, 38, 38, 33, 41, 42, 42, 41, 45, 45, 32, 48, 49, 50, 50, 49, 53, 53, 48, 56, 57, 57, 56, 60, 60),
                (-1, 0, 1, 2, 3, 4, 4, 3, 7, 7, 2, 10, 11, 11, 10, 14, 14, 1, 17, 18, 19, 19, 18, 22, 22, 17, 25, 26, 26, 25, 29, 29, 0, 32, 33, 34, 35, 35, 34, 38, 38, 33, 41, 42, 42, 41, 45, 45, 32, 48, 49, 50, 50, 49, 53, 53, 48, 56, 57, 57, 56, 60, 60)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 1, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5),
                (0, 1, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 1, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5),
                (0, 1, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 1, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5, 2, 3, 4, 5, 5, 4, 5, 5, 3, 4, 5, 5, 4, 5, 5)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((5, 6, 8, 9, 12, 13, 15, 16, 20, 21, 23, 24, 27, 28, 30, 31, 36, 37, 39, 40, 43, 44, 46, 47, 51, 52, 54, 55, 58, 59, 61, 62),
                (5, 6, 8, 9, 12, 13, 15, 16, 20, 21, 23, 24, 27, 28, 30, 31, 36, 37, 39, 40, 43, 44, 46, 47, 51, 52, 54, 55, 58, 59, 61, 62),
                (5, 6, 8, 9, 12, 13, 15, 16, 20, 21, 23, 24, 27, 28, 30, 31, 36, 37, 39, 40, 43, 44, 46, 47, 51, 52, 54, 55, 58, 59, 61, 62)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;